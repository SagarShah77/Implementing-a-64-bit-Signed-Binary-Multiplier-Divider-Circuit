
module muldiv ( result, valid, clock, reset, start, opera1, opera2, muordi );
  output [63:0] result;
  input [31:0] opera1;
  input [63:0] opera2;
  input clock, reset, start, muordi;
  output valid;
  wire   w4, \cust[1] , N145, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n259, n260, n284, n327, n329, n332, n335,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         \intadd_0/B[26] , \intadd_0/B[24] , \intadd_0/B[22] ,
         \intadd_0/B[20] , \intadd_0/B[18] , \intadd_0/B[16] ,
         \intadd_0/B[14] , \intadd_0/B[12] , \intadd_0/B[10] , \intadd_0/B[8] ,
         \intadd_0/B[6] , \intadd_0/B[4] , \intadd_0/B[2] , \intadd_0/B[0] ,
         \intadd_0/CI , \intadd_0/SUM[29] , \intadd_0/SUM[28] ,
         \intadd_0/SUM[27] , \intadd_0/SUM[26] , \intadd_0/SUM[25] ,
         \intadd_0/SUM[24] , \intadd_0/SUM[23] , \intadd_0/SUM[22] ,
         \intadd_0/SUM[21] , \intadd_0/SUM[20] , \intadd_0/SUM[19] ,
         \intadd_0/SUM[18] , \intadd_0/SUM[17] , \intadd_0/SUM[16] ,
         \intadd_0/SUM[15] , \intadd_0/SUM[14] , \intadd_0/SUM[13] ,
         \intadd_0/SUM[12] , \intadd_0/SUM[11] , \intadd_0/SUM[10] ,
         \intadd_0/SUM[9] , \intadd_0/SUM[8] , \intadd_0/SUM[7] ,
         \intadd_0/SUM[6] , \intadd_0/SUM[5] , \intadd_0/SUM[4] ,
         \intadd_0/SUM[3] , \intadd_0/SUM[2] , \intadd_0/SUM[1] ,
         \intadd_0/SUM[0] , \intadd_0/n30 , \intadd_0/n29 , \intadd_0/n28 ,
         \intadd_0/n27 , \intadd_0/n26 , \intadd_0/n25 , \intadd_0/n24 ,
         \intadd_0/n23 , \intadd_0/n22 , \intadd_0/n21 , \intadd_0/n20 ,
         \intadd_0/n19 , \intadd_0/n18 , \intadd_0/n17 , \intadd_0/n16 ,
         \intadd_0/n15 , \intadd_0/n14 , \intadd_0/n13 , \intadd_0/n12 ,
         \intadd_0/n11 , \intadd_0/n10 , \intadd_0/n9 , \intadd_0/n8 ,
         \intadd_0/n7 , \intadd_0/n6 , \intadd_0/n5 , \intadd_0/n4 ,
         \intadd_0/n3 , \intadd_0/n2 , \intadd_0/n1 , \intadd_1/CI ,
         \intadd_1/SUM[29] , \intadd_1/SUM[28] , \intadd_1/SUM[27] ,
         \intadd_1/SUM[26] , \intadd_1/SUM[25] , \intadd_1/SUM[24] ,
         \intadd_1/SUM[23] , \intadd_1/SUM[22] , \intadd_1/SUM[21] ,
         \intadd_1/SUM[20] , \intadd_1/SUM[19] , \intadd_1/SUM[18] ,
         \intadd_1/SUM[17] , \intadd_1/SUM[16] , \intadd_1/SUM[15] ,
         \intadd_1/SUM[14] , \intadd_1/SUM[13] , \intadd_1/SUM[12] ,
         \intadd_1/SUM[11] , \intadd_1/SUM[10] , \intadd_1/SUM[9] ,
         \intadd_1/SUM[8] , \intadd_1/SUM[7] , \intadd_1/SUM[6] ,
         \intadd_1/SUM[5] , \intadd_1/SUM[4] , \intadd_1/SUM[3] ,
         \intadd_1/SUM[2] , \intadd_1/SUM[1] , \intadd_1/SUM[0] ,
         \intadd_1/n30 , \intadd_1/n29 , \intadd_1/n28 , \intadd_1/n27 ,
         \intadd_1/n26 , \intadd_1/n25 , \intadd_1/n24 , \intadd_1/n23 ,
         \intadd_1/n22 , \intadd_1/n21 , \intadd_1/n20 , \intadd_1/n19 ,
         \intadd_1/n18 , \intadd_1/n17 , \intadd_1/n16 , \intadd_1/n15 ,
         \intadd_1/n14 , \intadd_1/n13 , \intadd_1/n12 , \intadd_1/n11 ,
         \intadd_1/n10 , \intadd_1/n9 , \intadd_1/n8 , \intadd_1/n7 ,
         \intadd_1/n6 , \intadd_1/n5 , \intadd_1/n4 , \intadd_1/n3 ,
         \intadd_1/n2 , \intadd_1/n1 , n1734, n1741, n1770, n1772, n1773,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n3076, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3275, n3276, n3277, n3278,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3956, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192;
  wire   [63:0] result_not;
  wire   [2:0] nest;
  wire   [31:0] D;
  wire   [31:0] result_copy;
  wire   [31:0] i;
  wire   [31:0] opera1_copy;
  wire   [31:0] opera1_copydiv;
  tri   cin1a;
  tri   cin1b;
  tri   cin2a;
  tri   cina;

  CTSX2 A8 ( .A(1'b0), .E(n3475), .Z(cina) );
  CTSX2 A7 ( .A(1'b1), .E(w4), .Z(cina) );
  CTSX2 A4 ( .A(1'b0), .E(n4986), .Z(cin1b) );
  CTSX2 A3 ( .A(1'b1), .E(n3136), .Z(cin1b) );
  CTSX2 A6 ( .A(1'b0), .E(n4478), .Z(cin2a) );
  CTSX2 A5 ( .A(1'b1), .E(n4479), .Z(cin2a) );
  CTSX2 A2 ( .A(1'b0), .E(n3136), .Z(cin1a) );
  CTSX2 A1 ( .A(1'b1), .E(n4986), .Z(cin1a) );
  CFA1X1 \intadd_0/U30  ( .A(n3468), .B(\intadd_0/n30 ), .CI(n3477), .CO(
        \intadd_0/n29 ), .S(\intadd_0/SUM[1] ) );
  CFA1X1 \intadd_0/U28  ( .A(n3469), .B(\intadd_0/n28 ), .CI(n1741), .CO(
        \intadd_0/n27 ), .S(\intadd_0/SUM[3] ) );
  CFA1X1 \intadd_0/U26  ( .A(n3456), .B(\intadd_0/n26 ), .CI(n3478), .CO(
        \intadd_0/n25 ), .S(\intadd_0/SUM[5] ) );
  CFA1X1 \intadd_0/U24  ( .A(n3457), .B(\intadd_0/n24 ), .CI(n3466), .CO(
        \intadd_0/n23 ), .S(\intadd_0/SUM[7] ) );
  CFA1X1 \intadd_0/U22  ( .A(n3458), .B(\intadd_0/n22 ), .CI(n3465), .CO(
        \intadd_0/n21 ), .S(\intadd_0/SUM[9] ) );
  CFA1X1 \intadd_0/U20  ( .A(n3459), .B(\intadd_0/n20 ), .CI(n3464), .CO(
        \intadd_0/n19 ), .S(\intadd_0/SUM[11] ) );
  CFA1X1 \intadd_0/U18  ( .A(n3443), .B(\intadd_0/n18 ), .CI(n3453), .CO(
        \intadd_0/n17 ), .S(\intadd_0/SUM[13] ) );
  CFA1X1 \intadd_0/U16  ( .A(n3444), .B(\intadd_0/n16 ), .CI(n3452), .CO(
        \intadd_0/n15 ), .S(\intadd_0/SUM[15] ) );
  CFA1X1 \intadd_0/U14  ( .A(n3445), .B(\intadd_0/n14 ), .CI(n3451), .CO(
        \intadd_0/n13 ), .S(\intadd_0/SUM[17] ) );
  CFA1X1 \intadd_0/U12  ( .A(n3399), .B(\intadd_0/n12 ), .CI(n3426), .CO(
        \intadd_0/n11 ), .S(\intadd_0/SUM[19] ) );
  CFA1X1 \intadd_0/U10  ( .A(n3400), .B(\intadd_0/n10 ), .CI(n3424), .CO(
        \intadd_0/n9 ), .S(\intadd_0/SUM[21] ) );
  CFA1X1 \intadd_0/U8  ( .A(n3401), .B(\intadd_0/n8 ), .CI(n3423), .CO(
        \intadd_0/n7 ), .S(\intadd_0/SUM[23] ) );
  CFA1X1 \intadd_0/U6  ( .A(n3383), .B(\intadd_0/n6 ), .CI(n3392), .CO(
        \intadd_0/n5 ), .S(\intadd_0/SUM[25] ) );
  CFA1X1 \intadd_0/U4  ( .A(n3384), .B(\intadd_0/n4 ), .CI(n3391), .CO(
        \intadd_0/n3 ), .S(\intadd_0/SUM[27] ) );
  CFA1X1 \intadd_0/U2  ( .A(n3385), .B(\intadd_0/n2 ), .CI(n3393), .CO(
        \intadd_0/n1 ), .S(\intadd_0/SUM[29] ) );
  CFA1X1 \intadd_1/U31  ( .A(n3316), .B(\intadd_1/CI ), .CI(n3473), .CO(
        \intadd_1/n30 ), .S(\intadd_1/SUM[0] ) );
  CFA1X1 \intadd_1/U30  ( .A(n3477), .B(\intadd_1/n30 ), .CI(n3467), .CO(
        \intadd_1/n29 ), .S(\intadd_1/SUM[1] ) );
  CFA1X1 \intadd_1/U29  ( .A(n3272), .B(\intadd_1/n29 ), .CI(n3472), .CO(
        \intadd_1/n28 ), .S(\intadd_1/SUM[2] ) );
  CFA1X1 \intadd_1/U28  ( .A(n1741), .B(\intadd_1/n28 ), .CI(n3471), .CO(
        \intadd_1/n27 ), .S(\intadd_1/SUM[3] ) );
  CFA1X1 \intadd_1/U27  ( .A(n3266), .B(\intadd_1/n27 ), .CI(n3470), .CO(
        \intadd_1/n26 ), .S(\intadd_1/SUM[4] ) );
  CFA1X1 \intadd_1/U26  ( .A(n3478), .B(\intadd_1/n26 ), .CI(n3455), .CO(
        \intadd_1/n25 ), .S(\intadd_1/SUM[5] ) );
  CFA1X1 \intadd_1/U25  ( .A(n3261), .B(\intadd_1/n25 ), .CI(n3463), .CO(
        \intadd_1/n24 ), .S(\intadd_1/SUM[6] ) );
  CFA1X1 \intadd_1/U24  ( .A(n3466), .B(\intadd_1/n24 ), .CI(n3462), .CO(
        \intadd_1/n23 ), .S(\intadd_1/SUM[7] ) );
  CFA1X1 \intadd_1/U23  ( .A(n3256), .B(\intadd_1/n23 ), .CI(n3460), .CO(
        \intadd_1/n22 ), .S(\intadd_1/SUM[8] ) );
  CFA1X1 \intadd_1/U22  ( .A(n3465), .B(\intadd_1/n22 ), .CI(n3454), .CO(
        \intadd_1/n21 ), .S(\intadd_1/SUM[9] ) );
  CFA1X1 \intadd_1/U21  ( .A(n3251), .B(\intadd_1/n21 ), .CI(n3461), .CO(
        \intadd_1/n20 ), .S(\intadd_1/SUM[10] ) );
  CFA1X1 \intadd_1/U20  ( .A(n3464), .B(\intadd_1/n20 ), .CI(n3450), .CO(
        \intadd_1/n19 ), .S(\intadd_1/SUM[11] ) );
  CFA1X1 \intadd_1/U19  ( .A(n3246), .B(\intadd_1/n19 ), .CI(n3447), .CO(
        \intadd_1/n18 ), .S(\intadd_1/SUM[12] ) );
  CFA1X1 \intadd_1/U18  ( .A(n3453), .B(\intadd_1/n18 ), .CI(n3442), .CO(
        \intadd_1/n17 ), .S(\intadd_1/SUM[13] ) );
  CFA1X1 \intadd_1/U17  ( .A(n3241), .B(\intadd_1/n17 ), .CI(n3449), .CO(
        \intadd_1/n16 ), .S(\intadd_1/SUM[14] ) );
  CFA1X1 \intadd_1/U16  ( .A(n3452), .B(\intadd_1/n16 ), .CI(n3448), .CO(
        \intadd_1/n15 ), .S(\intadd_1/SUM[15] ) );
  CFA1X1 \intadd_1/U15  ( .A(n3236), .B(\intadd_1/n15 ), .CI(n3446), .CO(
        \intadd_1/n14 ), .S(\intadd_1/SUM[16] ) );
  CFA1X1 \intadd_1/U14  ( .A(n3451), .B(\intadd_1/n14 ), .CI(n3441), .CO(
        \intadd_1/n13 ), .S(\intadd_1/SUM[17] ) );
  CFA1X1 \intadd_1/U13  ( .A(n3231), .B(\intadd_1/n13 ), .CI(n3406), .CO(
        \intadd_1/n12 ), .S(\intadd_1/SUM[18] ) );
  CFA1X1 \intadd_1/U12  ( .A(n3426), .B(\intadd_1/n12 ), .CI(n3405), .CO(
        \intadd_1/n11 ), .S(\intadd_1/SUM[19] ) );
  CFA1X1 \intadd_1/U11  ( .A(n3226), .B(\intadd_1/n11 ), .CI(n3402), .CO(
        \intadd_1/n10 ), .S(\intadd_1/SUM[20] ) );
  CFA1X1 \intadd_1/U10  ( .A(n3424), .B(\intadd_1/n10 ), .CI(n3398), .CO(
        \intadd_1/n9 ), .S(\intadd_1/SUM[21] ) );
  CFA1X1 \intadd_1/U9  ( .A(n3221), .B(\intadd_1/n9 ), .CI(n3404), .CO(
        \intadd_1/n8 ), .S(\intadd_1/SUM[22] ) );
  CFA1X1 \intadd_1/U8  ( .A(n3423), .B(\intadd_1/n8 ), .CI(n3403), .CO(
        \intadd_1/n7 ), .S(\intadd_1/SUM[23] ) );
  CFA1X1 \intadd_1/U7  ( .A(n3216), .B(\intadd_1/n7 ), .CI(n3386), .CO(
        \intadd_1/n6 ), .S(\intadd_1/SUM[24] ) );
  CFA1X1 \intadd_1/U6  ( .A(n3392), .B(\intadd_1/n6 ), .CI(n3382), .CO(
        \intadd_1/n5 ), .S(\intadd_1/SUM[25] ) );
  CFA1X1 \intadd_1/U5  ( .A(n3211), .B(\intadd_1/n5 ), .CI(n3388), .CO(
        \intadd_1/n4 ), .S(\intadd_1/SUM[26] ) );
  CFA1X1 \intadd_1/U4  ( .A(n3391), .B(\intadd_1/n4 ), .CI(n3381), .CO(
        \intadd_1/n3 ), .S(\intadd_1/SUM[27] ) );
  CFA1X1 \intadd_1/U3  ( .A(n3397), .B(\intadd_1/n3 ), .CI(n3387), .CO(
        \intadd_1/n2 ), .S(\intadd_1/SUM[28] ) );
  CFA1X1 \intadd_1/U2  ( .A(n3380), .B(\intadd_1/n2 ), .CI(n3393), .CO(
        \intadd_1/n1 ), .S(\intadd_1/SUM[29] ) );
  CFA1X1 \intadd_0/U31  ( .A(\intadd_0/B[0] ), .B(\intadd_0/CI ), .CI(n3316), 
        .CO(\intadd_0/n30 ), .S(\intadd_0/SUM[0] ) );
  CFA1X1 \intadd_0/U29  ( .A(\intadd_0/B[2] ), .B(\intadd_0/n29 ), .CI(n3272), 
        .CO(\intadd_0/n28 ), .S(\intadd_0/SUM[2] ) );
  CFA1X1 \intadd_0/U27  ( .A(\intadd_0/B[4] ), .B(\intadd_0/n27 ), .CI(n3266), 
        .CO(\intadd_0/n26 ), .S(\intadd_0/SUM[4] ) );
  CFA1X1 \intadd_0/U25  ( .A(\intadd_0/B[6] ), .B(\intadd_0/n25 ), .CI(n3261), 
        .CO(\intadd_0/n24 ), .S(\intadd_0/SUM[6] ) );
  CFA1X1 \intadd_0/U23  ( .A(\intadd_0/B[8] ), .B(\intadd_0/n23 ), .CI(n3256), 
        .CO(\intadd_0/n22 ), .S(\intadd_0/SUM[8] ) );
  CFA1X1 \intadd_0/U21  ( .A(\intadd_0/B[10] ), .B(\intadd_0/n21 ), .CI(n3251), 
        .CO(\intadd_0/n20 ), .S(\intadd_0/SUM[10] ) );
  CFA1X1 \intadd_0/U19  ( .A(\intadd_0/B[12] ), .B(\intadd_0/n19 ), .CI(n3246), 
        .CO(\intadd_0/n18 ), .S(\intadd_0/SUM[12] ) );
  CFA1X1 \intadd_0/U17  ( .A(\intadd_0/B[14] ), .B(\intadd_0/n17 ), .CI(n3241), 
        .CO(\intadd_0/n16 ), .S(\intadd_0/SUM[14] ) );
  CFA1X1 \intadd_0/U15  ( .A(\intadd_0/B[16] ), .B(\intadd_0/n15 ), .CI(n3236), 
        .CO(\intadd_0/n14 ), .S(\intadd_0/SUM[16] ) );
  CFA1X1 \intadd_0/U13  ( .A(\intadd_0/B[18] ), .B(\intadd_0/n13 ), .CI(n3231), 
        .CO(\intadd_0/n12 ), .S(\intadd_0/SUM[18] ) );
  CFA1X1 \intadd_0/U11  ( .A(\intadd_0/B[20] ), .B(\intadd_0/n11 ), .CI(n3226), 
        .CO(\intadd_0/n10 ), .S(\intadd_0/SUM[20] ) );
  CFA1X1 \intadd_0/U9  ( .A(\intadd_0/B[22] ), .B(\intadd_0/n9 ), .CI(n3221), 
        .CO(\intadd_0/n8 ), .S(\intadd_0/SUM[22] ) );
  CFA1X1 \intadd_0/U7  ( .A(\intadd_0/B[24] ), .B(\intadd_0/n7 ), .CI(n3216), 
        .CO(\intadd_0/n6 ), .S(\intadd_0/SUM[24] ) );
  CFA1X1 \intadd_0/U5  ( .A(\intadd_0/B[26] ), .B(\intadd_0/n5 ), .CI(n3211), 
        .CO(\intadd_0/n4 ), .S(\intadd_0/SUM[26] ) );
  CFA1X1 \intadd_0/U3  ( .A(n1772), .B(\intadd_0/n3 ), .CI(n3397), .CO(
        \intadd_0/n2 ), .S(\intadd_0/SUM[28] ) );
  CIVX2 U2842 ( .A(reset), .Z(n3076) );
  CIVX2 U2844 ( .A(n4468), .Z(n3078) );
  CIVX2 U2845 ( .A(n4169), .Z(n3079) );
  CIVX2 U2846 ( .A(n3648), .Z(n3080) );
  CIVX2 U2847 ( .A(n3738), .Z(n3081) );
  CIVX2 U2848 ( .A(n3743), .Z(n3082) );
  CIVX2 U2849 ( .A(n3749), .Z(n3083) );
  CIVX2 U2850 ( .A(n3497), .Z(n3084) );
  CIVX2 U2851 ( .A(n3487), .Z(n3085) );
  CIVX2 U2852 ( .A(n3599), .Z(n3086) );
  CIVX2 U2853 ( .A(n3579), .Z(n3087) );
  CIVX2 U2854 ( .A(n3559), .Z(n3088) );
  CIVX2 U2855 ( .A(n3538), .Z(n3089) );
  CIVX2 U2856 ( .A(n3501), .Z(n3090) );
  CIVX2 U2857 ( .A(n3513), .Z(n3091) );
  CIVX2 U2858 ( .A(n3523), .Z(n3092) );
  CIVX2 U2859 ( .A(n3533), .Z(n3093) );
  CIVX2 U2860 ( .A(n3544), .Z(n3094) );
  CIVX2 U2861 ( .A(n3556), .Z(n3095) );
  CIVX2 U2862 ( .A(n3565), .Z(n3096) );
  CIVX2 U2863 ( .A(n3576), .Z(n3097) );
  CIVX2 U2864 ( .A(n3585), .Z(n3098) );
  CIVX2 U2865 ( .A(n3596), .Z(n3099) );
  CIVX2 U2866 ( .A(n3619), .Z(n3100) );
  CIVX2 U2867 ( .A(n3605), .Z(n3101) );
  CIVX2 U2868 ( .A(n3616), .Z(n3102) );
  CIVX2 U2871 ( .A(n3733), .Z(n3105) );
  CIVX2 U2872 ( .A(n3727), .Z(n3106) );
  CIVX2 U2873 ( .A(n3724), .Z(n3107) );
  CIVX2 U2874 ( .A(n3721), .Z(n3108) );
  CIVX2 U2875 ( .A(n3718), .Z(n3109) );
  CIVX2 U2876 ( .A(n3715), .Z(n3110) );
  CIVX2 U2877 ( .A(n3710), .Z(n3111) );
  CIVX2 U2878 ( .A(n3707), .Z(n3112) );
  CIVX2 U2879 ( .A(n3704), .Z(n3113) );
  CIVX2 U2880 ( .A(n3699), .Z(n3114) );
  CIVX2 U2881 ( .A(n3696), .Z(n3115) );
  CIVX2 U2882 ( .A(n3693), .Z(n3116) );
  CIVX2 U2883 ( .A(n3688), .Z(n3117) );
  CIVX2 U2884 ( .A(n3685), .Z(n3118) );
  CIVX2 U2885 ( .A(n3682), .Z(n3119) );
  CIVX2 U2886 ( .A(n3677), .Z(n3120) );
  CIVX2 U2887 ( .A(n3674), .Z(n3121) );
  CIVX2 U2888 ( .A(n3671), .Z(n3122) );
  CIVX2 U2889 ( .A(n3666), .Z(n3123) );
  CIVX2 U2890 ( .A(n3663), .Z(n3124) );
  CIVX2 U2891 ( .A(n3660), .Z(n3125) );
  CIVX2 U2892 ( .A(n3625), .Z(n3126) );
  CIVX2 U2893 ( .A(n3492), .Z(n3127) );
  CIVX2 U2895 ( .A(n3655), .Z(n3129) );
  CIVX2 U2896 ( .A(n3650), .Z(n3130) );
  CIVX2 U2897 ( .A(n3635), .Z(n3131) );
  CIVX2 U2898 ( .A(n3652), .Z(n3132) );
  CIVX2 U2899 ( .A(n3668), .Z(n3133) );
  CIVX2 U2900 ( .A(n3690), .Z(n3134) );
  CIVX2 U2901 ( .A(n3712), .Z(n3135) );
  CIVX2 U2902 ( .A(n4986), .Z(n3136) );
  CIVX2 U2903 ( .A(n4690), .Z(n3137) );
  CIVX2 U2904 ( .A(n4694), .Z(n3138) );
  CIVX2 U2905 ( .A(n4571), .Z(n3139) );
  CIVX2 U2906 ( .A(n4700), .Z(n3140) );
  CIVX2 U2907 ( .A(n4568), .Z(n3141) );
  CIVX2 U2908 ( .A(n4812), .Z(n3142) );
  CIVX2 U2909 ( .A(n4728), .Z(n3143) );
  CIVX2 U2910 ( .A(n4818), .Z(n3144) );
  CIVX2 U2911 ( .A(n4720), .Z(n3145) );
  CIVX2 U2912 ( .A(n4817), .Z(n3146) );
  CIVX2 U2913 ( .A(n4734), .Z(n3147) );
  CIVX2 U2914 ( .A(n4870), .Z(n3148) );
  CIVX2 U2915 ( .A(n4841), .Z(n3149) );
  CIVX2 U2916 ( .A(n4868), .Z(n3150) );
  CIVX2 U2917 ( .A(n4865), .Z(n3151) );
  CIVX2 U2918 ( .A(n4875), .Z(n3152) );
  CIVX2 U2919 ( .A(n4836), .Z(n3153) );
  CIVX2 U2920 ( .A(n4863), .Z(n3154) );
  CIVX2 U2921 ( .A(n4899), .Z(n3155) );
  CIVX2 U2922 ( .A(n4928), .Z(n3156) );
  CIVX2 U2923 ( .A(n4895), .Z(n3157) );
  CIVX2 U2924 ( .A(n4921), .Z(n3158) );
  CIVX2 U2925 ( .A(n4923), .Z(n3159) );
  CIVX2 U2926 ( .A(n4935), .Z(n3160) );
  CIVX2 U2927 ( .A(n4969), .Z(n3161) );
  CIVX2 U2928 ( .A(n4977), .Z(n3162) );
  CIVX2 U2929 ( .A(n4943), .Z(n3163) );
  CIVX2 U2930 ( .A(n4971), .Z(n3164) );
  CIVX2 U2932 ( .A(n3773), .Z(n3166) );
  CIVX2 U2933 ( .A(n3947), .Z(n3167) );
  CIVX2 U2934 ( .A(n3920), .Z(n3168) );
  CIVX2 U2935 ( .A(n3909), .Z(n3169) );
  CIVX2 U2936 ( .A(n3899), .Z(n3170) );
  CIVX2 U2937 ( .A(n3888), .Z(n3171) );
  CIVX2 U2938 ( .A(n3878), .Z(n3172) );
  CIVX2 U2939 ( .A(n3867), .Z(n3173) );
  CIVX2 U2940 ( .A(n3857), .Z(n3174) );
  CIVX2 U2941 ( .A(n3846), .Z(n3175) );
  CIVX2 U2942 ( .A(n3836), .Z(n3176) );
  CIVX2 U2943 ( .A(n3819), .Z(n3177) );
  CIVX2 U2944 ( .A(n3777), .Z(n3178) );
  CIVX2 U2945 ( .A(n3780), .Z(n3179) );
  CIVX2 U2947 ( .A(n5096), .Z(n3181) );
  CIVX2 U2948 ( .A(n5090), .Z(n3182) );
  CIVX2 U2949 ( .A(n5085), .Z(n3183) );
  CIVX2 U2950 ( .A(n4507), .Z(n3184) );
  CIVX2 U2951 ( .A(n5079), .Z(n3185) );
  CIVX2 U2952 ( .A(n4517), .Z(n3186) );
  CIVX2 U2953 ( .A(n4515), .Z(n3187) );
  CIVX2 U2954 ( .A(n5068), .Z(n3188) );
  CIVX2 U2955 ( .A(n4513), .Z(n3189) );
  CIVX2 U2956 ( .A(n4505), .Z(n3190) );
  CIVX2 U2957 ( .A(n5058), .Z(n3191) );
  CIVX2 U2958 ( .A(n4511), .Z(n3192) );
  CIVX2 U2959 ( .A(n4503), .Z(n3193) );
  CIVX2 U2960 ( .A(n4539), .Z(n3194) );
  CIVX2 U2961 ( .A(n4521), .Z(n3195) );
  CIVX2 U2962 ( .A(n5040), .Z(n3196) );
  CIVX2 U2963 ( .A(n4526), .Z(n3197) );
  CIVX2 U2964 ( .A(n4708), .Z(n3198) );
  CIVX2 U2967 ( .A(n3763), .Z(n3201) );
  CIVX2 U2968 ( .A(\intadd_0/SUM[29] ), .Z(n3202) );
  CIVX2 U2969 ( .A(\intadd_0/SUM[28] ), .Z(n3203) );
  CIVX2 U2970 ( .A(\intadd_0/SUM[27] ), .Z(n3204) );
  CIVX2 U2971 ( .A(\intadd_0/SUM[26] ), .Z(n3205) );
  CIVX2 U2972 ( .A(n3759), .Z(n3206) );
  CIVX2 U2973 ( .A(\intadd_1/SUM[29] ), .Z(n3207) );
  CIVX2 U2974 ( .A(\intadd_1/SUM[28] ), .Z(n3208) );
  CIVX2 U2975 ( .A(\intadd_1/SUM[27] ), .Z(n3209) );
  CIVX2 U2976 ( .A(\intadd_1/SUM[26] ), .Z(n3210) );
  CIVX2 U2978 ( .A(\intadd_0/SUM[25] ), .Z(n3212) );
  CIVX2 U2979 ( .A(\intadd_0/SUM[24] ), .Z(n3213) );
  CIVX2 U2980 ( .A(\intadd_1/SUM[25] ), .Z(n3214) );
  CIVX2 U2981 ( .A(\intadd_1/SUM[24] ), .Z(n3215) );
  CIVX2 U2983 ( .A(\intadd_0/SUM[23] ), .Z(n3217) );
  CIVX2 U2984 ( .A(\intadd_0/SUM[22] ), .Z(n3218) );
  CIVX2 U2985 ( .A(\intadd_1/SUM[23] ), .Z(n3219) );
  CIVX2 U2986 ( .A(\intadd_1/SUM[22] ), .Z(n3220) );
  CIVX2 U2988 ( .A(\intadd_0/SUM[21] ), .Z(n3222) );
  CIVX2 U2989 ( .A(\intadd_0/SUM[20] ), .Z(n3223) );
  CIVX2 U2990 ( .A(\intadd_1/SUM[21] ), .Z(n3224) );
  CIVX2 U2991 ( .A(\intadd_1/SUM[20] ), .Z(n3225) );
  CIVX2 U2993 ( .A(\intadd_0/SUM[19] ), .Z(n3227) );
  CIVX2 U2994 ( .A(\intadd_0/SUM[18] ), .Z(n3228) );
  CIVX2 U2995 ( .A(\intadd_1/SUM[19] ), .Z(n3229) );
  CIVX2 U2996 ( .A(\intadd_1/SUM[18] ), .Z(n3230) );
  CIVX2 U2998 ( .A(\intadd_0/SUM[17] ), .Z(n3232) );
  CIVX2 U2999 ( .A(\intadd_0/SUM[16] ), .Z(n3233) );
  CIVX2 U3000 ( .A(\intadd_1/SUM[17] ), .Z(n3234) );
  CIVX2 U3001 ( .A(\intadd_1/SUM[16] ), .Z(n3235) );
  CIVX2 U3003 ( .A(\intadd_0/SUM[15] ), .Z(n3237) );
  CIVX2 U3004 ( .A(\intadd_0/SUM[14] ), .Z(n3238) );
  CIVX2 U3005 ( .A(\intadd_1/SUM[15] ), .Z(n3239) );
  CIVX2 U3006 ( .A(\intadd_1/SUM[14] ), .Z(n3240) );
  CIVX2 U3008 ( .A(\intadd_0/SUM[13] ), .Z(n3242) );
  CIVX2 U3009 ( .A(\intadd_0/SUM[12] ), .Z(n3243) );
  CIVX2 U3010 ( .A(\intadd_1/SUM[13] ), .Z(n3244) );
  CIVX2 U3011 ( .A(\intadd_1/SUM[12] ), .Z(n3245) );
  CIVX2 U3013 ( .A(\intadd_0/SUM[11] ), .Z(n3247) );
  CIVX2 U3014 ( .A(\intadd_0/SUM[10] ), .Z(n3248) );
  CIVX2 U3015 ( .A(\intadd_1/SUM[11] ), .Z(n3249) );
  CIVX2 U3016 ( .A(\intadd_1/SUM[10] ), .Z(n3250) );
  CIVX2 U3018 ( .A(\intadd_0/SUM[9] ), .Z(n3252) );
  CIVX2 U3019 ( .A(\intadd_0/SUM[8] ), .Z(n3253) );
  CIVX2 U3020 ( .A(\intadd_1/SUM[9] ), .Z(n3254) );
  CIVX2 U3021 ( .A(\intadd_1/SUM[8] ), .Z(n3255) );
  CIVX2 U3023 ( .A(\intadd_0/SUM[7] ), .Z(n3257) );
  CIVX2 U3024 ( .A(\intadd_0/SUM[6] ), .Z(n3258) );
  CIVX2 U3025 ( .A(\intadd_1/SUM[7] ), .Z(n3259) );
  CIVX2 U3026 ( .A(\intadd_1/SUM[6] ), .Z(n3260) );
  CIVX2 U3028 ( .A(\intadd_0/SUM[5] ), .Z(n3262) );
  CIVX2 U3029 ( .A(\intadd_0/SUM[4] ), .Z(n3263) );
  CIVX2 U3030 ( .A(\intadd_1/SUM[5] ), .Z(n3264) );
  CIVX2 U3031 ( .A(\intadd_1/SUM[4] ), .Z(n3265) );
  CIVX2 U3033 ( .A(\intadd_0/SUM[3] ), .Z(n3267) );
  CIVX2 U3034 ( .A(\intadd_0/SUM[2] ), .Z(n3268) );
  CIVX2 U3035 ( .A(\intadd_1/SUM[3] ), .Z(n3269) );
  CIVX2 U3036 ( .A(\intadd_1/SUM[2] ), .Z(n3270) );
  CIVX2 U3037 ( .A(n3973), .Z(n3271) );
  CIVX2 U3041 ( .A(n3949), .Z(n3275) );
  CIVX2 U3043 ( .A(n3967), .Z(n3277) );
  CIVX2 U3044 ( .A(n3766), .Z(n3278) );
  CIVX2 U3049 ( .A(i[3]), .Z(n3283) );
  CIVX2 U3050 ( .A(n5009), .Z(n3284) );
  CIVX2 U3051 ( .A(result_copy[27]), .Z(n3285) );
  CIVX2 U3052 ( .A(result_copy[25]), .Z(n3286) );
  CIVX2 U3053 ( .A(result_copy[17]), .Z(n3287) );
  CIVX2 U3054 ( .A(result_copy[13]), .Z(n3288) );
  CIVX2 U3055 ( .A(result_copy[9]), .Z(n3289) );
  CIVX2 U3056 ( .A(result_copy[5]), .Z(n3290) );
  CIVX2 U3057 ( .A(result_copy[1]), .Z(n3291) );
  CIVX2 U3058 ( .A(n4462), .Z(n3292) );
  CIVX2 U3059 ( .A(result_copy[29]), .Z(n3293) );
  CIVX2 U3060 ( .A(result_copy[21]), .Z(n3294) );
  CIVX2 U3061 ( .A(result_copy[19]), .Z(n3295) );
  CIVX2 U3062 ( .A(result_copy[23]), .Z(n3296) );
  CIVX2 U3063 ( .A(n4469), .Z(n3297) );
  CIVX2 U3064 ( .A(n4459), .Z(n3298) );
  CIVX2 U3065 ( .A(n4456), .Z(n3299) );
  CIVX2 U3066 ( .A(n4453), .Z(n3300) );
  CIVX2 U3067 ( .A(n4450), .Z(n3301) );
  CIVX2 U3068 ( .A(n4447), .Z(n3302) );
  CIVX2 U3069 ( .A(n4444), .Z(n3303) );
  CIVX2 U3070 ( .A(n4441), .Z(n3304) );
  CIVX2 U3071 ( .A(n4438), .Z(n3305) );
  CIVX2 U3072 ( .A(n4435), .Z(n3306) );
  CIVX2 U3073 ( .A(n4432), .Z(n3307) );
  CIVX2 U3074 ( .A(n4429), .Z(n3308) );
  CIVX2 U3075 ( .A(n4426), .Z(n3309) );
  CIVX2 U3076 ( .A(n4423), .Z(n3310) );
  CIVX2 U3077 ( .A(n4420), .Z(n3311) );
  CIVX2 U3078 ( .A(\intadd_0/SUM[1] ), .Z(n3312) );
  CIVX2 U3079 ( .A(\intadd_0/SUM[0] ), .Z(n3313) );
  CIVX2 U3080 ( .A(\intadd_1/SUM[1] ), .Z(n3314) );
  CIVX2 U3081 ( .A(\intadd_1/SUM[0] ), .Z(n3315) );
  CIVX2 U3084 ( .A(n4417), .Z(n3318) );
  CIVX2 U3085 ( .A(n4414), .Z(n3319) );
  CIVX2 U3086 ( .A(n4411), .Z(n3320) );
  CIVX2 U3087 ( .A(n4408), .Z(n3321) );
  CIVX2 U3088 ( .A(n4405), .Z(n3322) );
  CIVX2 U3089 ( .A(n4402), .Z(n3323) );
  CIVX2 U3090 ( .A(n4399), .Z(n3324) );
  CIVX2 U3091 ( .A(n4396), .Z(n3325) );
  CIVX2 U3092 ( .A(n4393), .Z(n3326) );
  CIVX2 U3093 ( .A(n4390), .Z(n3327) );
  CIVX2 U3094 ( .A(n4387), .Z(n3328) );
  CIVX2 U3095 ( .A(n4384), .Z(n3329) );
  CIVX2 U3096 ( .A(n4381), .Z(n3330) );
  CIVX2 U3097 ( .A(n4378), .Z(n3331) );
  CIVX2 U3098 ( .A(n4375), .Z(n3332) );
  CIVX2 U3099 ( .A(n4372), .Z(n3333) );
  CIVX2 U3100 ( .A(n4369), .Z(n3334) );
  CIVX2 U3101 ( .A(n4366), .Z(n3335) );
  CIVX2 U3102 ( .A(n4363), .Z(n3336) );
  CIVX2 U3103 ( .A(n4360), .Z(n3337) );
  CIVX2 U3104 ( .A(n4357), .Z(n3338) );
  CIVX2 U3105 ( .A(n4354), .Z(n3339) );
  CIVX2 U3106 ( .A(n4351), .Z(n3340) );
  CIVX2 U3107 ( .A(n4348), .Z(n3341) );
  CIVX2 U3108 ( .A(n4345), .Z(n3342) );
  CIVX2 U3109 ( .A(n4342), .Z(n3343) );
  CIVX2 U3110 ( .A(n4339), .Z(n3344) );
  CIVX2 U3111 ( .A(n4336), .Z(n3345) );
  CIVX2 U3112 ( .A(n4333), .Z(n3346) );
  CIVX2 U3113 ( .A(n4330), .Z(n3347) );
  CIVX2 U3114 ( .A(n4327), .Z(n3348) );
  CIVX2 U3115 ( .A(n4324), .Z(n3349) );
  CIVX2 U3116 ( .A(n4321), .Z(n3350) );
  CIVX2 U3117 ( .A(n4318), .Z(n3351) );
  CIVX2 U3118 ( .A(n4315), .Z(n3352) );
  CIVX2 U3119 ( .A(n4312), .Z(n3353) );
  CIVX2 U3120 ( .A(n4308), .Z(n3354) );
  CIVX2 U3121 ( .A(n4305), .Z(n3355) );
  CIVX2 U3122 ( .A(n4300), .Z(n3356) );
  CIVX2 U3123 ( .A(n4295), .Z(n3357) );
  CIVX2 U3124 ( .A(n4290), .Z(n3358) );
  CIVX2 U3125 ( .A(n4285), .Z(n3359) );
  CIVX2 U3126 ( .A(n3744), .Z(n3360) );
  CIVX2 U3127 ( .A(i[0]), .Z(n3361) );
  CIVX2 U3129 ( .A(n5007), .Z(n3363) );
  CIVX2 U3130 ( .A(result_copy[3]), .Z(n3364) );
  CIVX2 U3131 ( .A(result_copy[7]), .Z(n3365) );
  CIVX2 U3134 ( .A(result_copy[26]), .Z(n3366) );
  CIVX2 U3135 ( .A(result_copy[12]), .Z(n3367) );
  CIVX2 U3136 ( .A(result_copy[16]), .Z(n3368) );
  CIVX2 U3137 ( .A(result_copy[24]), .Z(n3369) );
  CIVX2 U3138 ( .A(result_copy[10]), .Z(n3370) );
  CIVX2 U3139 ( .A(result_copy[14]), .Z(n3371) );
  CIVX2 U3140 ( .A(result_copy[18]), .Z(n3372) );
  CIVX2 U3141 ( .A(result_copy[30]), .Z(n3373) );
  CIVX2 U3142 ( .A(result_copy[20]), .Z(n3374) );
  CIVX2 U3143 ( .A(result_copy[22]), .Z(n3375) );
  CIVX2 U3144 ( .A(result_copy[28]), .Z(n3376) );
  CIVX2 U3146 ( .A(n332), .Z(n3378) );
  CIVX2 U3147 ( .A(n329), .Z(n3379) );
  CIVX2 U3148 ( .A(opera1_copy[30]), .Z(n3380) );
  CIVX2 U3149 ( .A(opera1_copy[28]), .Z(n3381) );
  CIVX2 U3150 ( .A(opera1_copy[26]), .Z(n3382) );
  CIVX2 U3153 ( .A(opera1_copydiv[30]), .Z(n3385) );
  CIVX2 U3154 ( .A(opera1_copy[25]), .Z(n3386) );
  CIVX2 U3155 ( .A(opera1_copy[29]), .Z(n3387) );
  CIVX2 U3156 ( .A(opera1_copy[27]), .Z(n3388) );
  CIVX2 U3158 ( .A(opera1_copy[31]), .Z(n3390) );
  CIVX2 U3159 ( .A(D[28]), .Z(n3391) );
  CIVX2 U3160 ( .A(D[26]), .Z(n3392) );
  CIVX2 U3161 ( .A(D[30]), .Z(n3393) );
  CIVX2 U3162 ( .A(n3944), .Z(n3394) );
  CIVX2 U3163 ( .A(i[27]), .Z(n3395) );
  CIVX2 U3164 ( .A(D[31]), .Z(n3396) );
  CIVX2 U3166 ( .A(opera1_copy[22]), .Z(n3398) );
  CIVX2 U3167 ( .A(opera1_copydiv[20]), .Z(n3399) );
  CIVX2 U3169 ( .A(opera1_copydiv[24]), .Z(n3401) );
  CIVX2 U3170 ( .A(opera1_copy[21]), .Z(n3402) );
  CIVX2 U3171 ( .A(opera1_copy[24]), .Z(n3403) );
  CIVX2 U3172 ( .A(opera1_copy[23]), .Z(n3404) );
  CIVX2 U3173 ( .A(opera1_copy[20]), .Z(n3405) );
  CIVX2 U3174 ( .A(opera1_copy[19]), .Z(n3406) );
  CIVX2 U3175 ( .A(i[30]), .Z(n3407) );
  CIVX2 U3176 ( .A(i[22]), .Z(n3408) );
  CIVX2 U3177 ( .A(i[14]), .Z(n3409) );
  CIVX2 U3178 ( .A(i[8]), .Z(n3410) );
  CIVX2 U3179 ( .A(i[6]), .Z(n3411) );
  CIVX2 U3180 ( .A(i[16]), .Z(n3412) );
  CIVX2 U3182 ( .A(n3752), .Z(n3414) );
  CIVX2 U3183 ( .A(n4170), .Z(n3415) );
  CIVX2 U3184 ( .A(i[18]), .Z(n3416) );
  CIVX2 U3185 ( .A(i[20]), .Z(n3417) );
  CIVX2 U3186 ( .A(i[28]), .Z(n3418) );
  CIVX2 U3187 ( .A(i[24]), .Z(n3419) );
  CIVX2 U3188 ( .A(i[26]), .Z(n3420) );
  CIVX2 U3189 ( .A(i[10]), .Z(n3421) );
  CIVX2 U3190 ( .A(i[12]), .Z(n3422) );
  CIVX2 U3191 ( .A(D[24]), .Z(n3423) );
  CIVX2 U3192 ( .A(D[22]), .Z(n3424) );
  CIVX2 U3193 ( .A(i[29]), .Z(n3425) );
  CIVX2 U3194 ( .A(D[20]), .Z(n3426) );
  CIVX2 U3195 ( .A(i[7]), .Z(n3427) );
  CIVX2 U3196 ( .A(i[17]), .Z(n3428) );
  CIVX2 U3197 ( .A(i[9]), .Z(n3429) );
  CIVX2 U3198 ( .A(i[25]), .Z(n3430) );
  CIVX2 U3199 ( .A(i[13]), .Z(n3431) );
  CIVX2 U3200 ( .A(i[23]), .Z(n3432) );
  CIVX2 U3201 ( .A(i[11]), .Z(n3433) );
  CIVX2 U3202 ( .A(i[15]), .Z(n3434) );
  CIVX2 U3203 ( .A(i[21]), .Z(n3435) );
  CIVX2 U3204 ( .A(i[19]), .Z(n3436) );
  CIVX2 U3205 ( .A(i[2]), .Z(n3437) );
  CIVX2 U3206 ( .A(i[4]), .Z(n3438) );
  CIVX2 U3207 ( .A(i[5]), .Z(n3439) );
  CIVX2 U3209 ( .A(opera1_copy[18]), .Z(n3441) );
  CIVX2 U3210 ( .A(opera1_copy[14]), .Z(n3442) );
  CIVX2 U3212 ( .A(opera1_copydiv[16]), .Z(n3444) );
  CIVX2 U3214 ( .A(opera1_copy[17]), .Z(n3446) );
  CIVX2 U3215 ( .A(opera1_copy[13]), .Z(n3447) );
  CIVX2 U3216 ( .A(opera1_copy[16]), .Z(n3448) );
  CIVX2 U3217 ( .A(opera1_copy[15]), .Z(n3449) );
  CIVX2 U3218 ( .A(opera1_copy[12]), .Z(n3450) );
  CIVX2 U3219 ( .A(D[18]), .Z(n3451) );
  CIVX2 U3220 ( .A(D[16]), .Z(n3452) );
  CIVX2 U3221 ( .A(D[14]), .Z(n3453) );
  CIVX2 U3222 ( .A(opera1_copy[10]), .Z(n3454) );
  CIVX2 U3223 ( .A(opera1_copy[6]), .Z(n3455) );
  CIVX2 U3225 ( .A(opera1_copydiv[8]), .Z(n3457) );
  CIVX2 U3227 ( .A(opera1_copydiv[12]), .Z(n3459) );
  CIVX2 U3228 ( .A(opera1_copy[9]), .Z(n3460) );
  CIVX2 U3229 ( .A(opera1_copy[11]), .Z(n3461) );
  CIVX2 U3230 ( .A(opera1_copy[8]), .Z(n3462) );
  CIVX2 U3231 ( .A(opera1_copy[7]), .Z(n3463) );
  CIVX2 U3232 ( .A(D[12]), .Z(n3464) );
  CIVX2 U3233 ( .A(D[10]), .Z(n3465) );
  CIVX2 U3234 ( .A(D[8]), .Z(n3466) );
  CIVX2 U3235 ( .A(opera1_copy[2]), .Z(n3467) );
  CIVX2 U3236 ( .A(opera1_copydiv[2]), .Z(n3468) );
  CIVX2 U3237 ( .A(opera1_copydiv[4]), .Z(n3469) );
  CIVX2 U3238 ( .A(opera1_copy[5]), .Z(n3470) );
  CIVX2 U3239 ( .A(opera1_copy[4]), .Z(n3471) );
  CIVX2 U3240 ( .A(opera1_copy[3]), .Z(n3472) );
  CIVX2 U3241 ( .A(opera1_copy[1]), .Z(n3473) );
  CIVX2 U3243 ( .A(w4), .Z(n3475) );
  CIVX2 U3244 ( .A(n3945), .Z(n3476) );
  CIVX2 U3245 ( .A(D[2]), .Z(n3477) );
  CIVX2 U3246 ( .A(D[6]), .Z(n3478) );
  CIVX2 U3248 ( .A(result_copy[6]), .Z(n3480) );
  CIVX2 U3249 ( .A(result_copy[2]), .Z(n3481) );
  CIVX2 U3250 ( .A(D[0]), .Z(n3482) );
  CND2IX1 U3252 ( .B(n4984), .A(n3131), .Z(n3641) );
  COR4X1 U3253 ( .A(n3440), .B(n3361), .C(n3081), .D(i[2]), .Z(n3737) );
  COR4X1 U3254 ( .A(n3438), .B(n3283), .C(n3360), .D(n3081), .Z(n3750) );
  COR4X1 U3255 ( .A(n5190), .B(n3756), .C(n4481), .D(n3757), .Z(n1622) );
  CAOR1X1 U3256 ( .A(n3786), .B(n5182), .C(n3791), .Z(n3789) );
  CAOR1X1 U3257 ( .A(n4478), .B(n5052), .C(n3849), .Z(n3842) );
  CAOR1X1 U3258 ( .A(n4478), .B(n5063), .C(n3870), .Z(n3863) );
  CAOR1X1 U3259 ( .A(n4478), .B(n5074), .C(n3891), .Z(n3884) );
  CAOR1X1 U3260 ( .A(n4478), .B(n5085), .C(n3912), .Z(n3905) );
  CAOR2X1 U3261 ( .A(n5101), .B(n5180), .C(n3936), .D(n5181), .Z(n3935) );
  COR4X1 U3262 ( .A(n3974), .B(n3975), .C(n3976), .D(n3977), .Z(n1584) );
  COR4X1 U3263 ( .A(n4000), .B(n4001), .C(n4002), .D(n4003), .Z(n1580) );
  COR4X1 U3264 ( .A(n4026), .B(n4027), .C(n4028), .D(n4029), .Z(n1576) );
  COR4X1 U3265 ( .A(n4052), .B(n4053), .C(n4054), .D(n4055), .Z(n1572) );
  COR4X1 U3266 ( .A(n4078), .B(n4079), .C(n4080), .D(n4081), .Z(n1568) );
  COR4X1 U3267 ( .A(n4104), .B(n4105), .C(n4106), .D(n4107), .Z(n1564) );
  COR4X1 U3268 ( .A(n4130), .B(n4131), .C(n4132), .D(n4133), .Z(n1560) );
  CND2IX1 U3269 ( .B(n4150), .A(n4482), .Z(n3772) );
  CAOR1X1 U3270 ( .A(n4478), .B(n5052), .C(n3192), .Z(n4159) );
  CAOR1X1 U3271 ( .A(n4478), .B(n5063), .C(n3189), .Z(n4157) );
  CAOR1X1 U3272 ( .A(n4478), .B(n5074), .C(n3186), .Z(n4155) );
  COAN1X1 U3274 ( .A(opera1_copydiv[0]), .B(D[0]), .C(\intadd_0/CI ), .Z(n3948) );
  CND2IX1 U3275 ( .B(n4148), .A(n3414), .Z(n4168) );
  CAN4X1 U3276 ( .A(n3438), .B(n3283), .C(n3437), .D(n3440), .Z(n4275) );
  CFD1QXL \nest_reg[1]  ( .D(n3079), .CP(clock), .Q(nest[1]) );
  CFD1QXL \nest_reg[2]  ( .D(n1555), .CP(clock), .Q(nest[2]) );
  CFD1QXL \nest_reg[0]  ( .D(n1687), .CP(clock), .Q(nest[0]) );
  CFD1QXL \result_not_reg[63]  ( .D(n4490), .CP(clock), .Q(result_not[63]) );
  CFD1QXL \result_copy_reg[3]  ( .D(n4492), .CP(clock), .Q(result_copy[3]) );
  CFD1QXL \result_copy_reg[7]  ( .D(n4497), .CP(clock), .Q(result_copy[7]) );
  CFD1QXL \result_copy_reg[26]  ( .D(n4502), .CP(clock), .Q(result_copy[26])
         );
  CFD1QXL \result_copy_reg[12]  ( .D(n4504), .CP(clock), .Q(result_copy[12])
         );
  CFD1QXL \result_copy_reg[16]  ( .D(n4506), .CP(clock), .Q(result_copy[16])
         );
  CFD1QXL \result_copy_reg[24]  ( .D(n4508), .CP(clock), .Q(result_copy[24])
         );
  CFD1QXL \result_copy_reg[10]  ( .D(n4510), .CP(clock), .Q(result_copy[10])
         );
  CFD1QXL \result_copy_reg[14]  ( .D(n4512), .CP(clock), .Q(result_copy[14])
         );
  CFD1QXL \result_copy_reg[18]  ( .D(n4514), .CP(clock), .Q(result_copy[18])
         );
  CFD1QXL \result_copy_reg[20]  ( .D(n4516), .CP(clock), .Q(result_copy[20])
         );
  CFD1QXL \result_copy_reg[22]  ( .D(n4518), .CP(clock), .Q(result_copy[22])
         );
  CFD1QXL \result_copy_reg[28]  ( .D(n4520), .CP(clock), .Q(result_copy[28])
         );
  CFD1QXL \result_copy_reg[6]  ( .D(n4522), .CP(clock), .Q(result_copy[6]) );
  CFD1QXL \result_copy_reg[2]  ( .D(n4523), .CP(clock), .Q(result_copy[2]) );
  CFD1QXL \result_not_reg[62]  ( .D(n4527), .CP(clock), .Q(result_not[62]) );
  CFD1QXL \result_copy_reg[30]  ( .D(n4529), .CP(clock), .Q(result_copy[30])
         );
  CFD1XL \result_copy_reg[4]  ( .D(n4531), .CP(clock), .QN(n332) );
  CFD1XL \result_copy_reg[8]  ( .D(n4535), .CP(clock), .QN(n329) );
  CFD1XL \result_copy_reg[11]  ( .D(n4540), .CP(clock), .QN(n327) );
  CFD1QXL \result_reg[9]  ( .D(n4541), .CP(clock), .Q(result[9]) );
  CFD1QXL \result_reg[7]  ( .D(n4543), .CP(clock), .Q(result[7]) );
  CFD1QXL \result_reg[5]  ( .D(n4545), .CP(clock), .Q(result[5]) );
  CFD1QXL \result_reg[3]  ( .D(n4547), .CP(clock), .Q(result[3]) );
  CFD1QXL \result_reg[1]  ( .D(n4549), .CP(clock), .Q(result[1]) );
  CFD1QXL \result_reg[6]  ( .D(n4551), .CP(clock), .Q(result[6]) );
  CFD1QXL \result_reg[2]  ( .D(n4553), .CP(clock), .Q(result[2]) );
  CFD1QXL \result_reg[0]  ( .D(n4555), .CP(clock), .Q(result[0]) );
  CFD1QXL \result_reg[63]  ( .D(n4557), .CP(clock), .Q(result[63]) );
  CFD1QXL \result_reg[8]  ( .D(n4559), .CP(clock), .Q(result[8]) );
  CFD1QXL \result_reg[4]  ( .D(n4561), .CP(clock), .Q(result[4]) );
  CFD1QXL \opera1_copy_reg[30]  ( .D(n4563), .CP(clock), .Q(opera1_copy[30])
         );
  CFD1QXL \opera1_copy_reg[28]  ( .D(n4564), .CP(clock), .Q(opera1_copy[28])
         );
  CFD1QXL \opera1_copy_reg[26]  ( .D(n4566), .CP(clock), .Q(opera1_copy[26])
         );
  CFD1QXL \opera1_copydiv_reg[26]  ( .D(n4570), .CP(clock), .Q(
        opera1_copydiv[26]) );
  CFD1QXL \opera1_copydiv_reg[28]  ( .D(n4573), .CP(clock), .Q(
        opera1_copydiv[28]) );
  CFD1QXL \opera1_copydiv_reg[30]  ( .D(n4574), .CP(clock), .Q(
        opera1_copydiv[30]) );
  CFD1QXL \opera1_copy_reg[27]  ( .D(n4576), .CP(clock), .Q(opera1_copy[27])
         );
  CFD1QXL \opera1_copy_reg[31]  ( .D(n4579), .CP(clock), .Q(opera1_copy[31])
         );
  CFD1QXL \result_reg[31]  ( .D(n4580), .CP(clock), .Q(result[31]) );
  CFD1QXL \result_reg[29]  ( .D(n4582), .CP(clock), .Q(result[29]) );
  CFD1QXL \result_reg[27]  ( .D(n4584), .CP(clock), .Q(result[27]) );
  CFD1QXL \result_reg[25]  ( .D(n4586), .CP(clock), .Q(result[25]) );
  CFD1QXL \result_reg[23]  ( .D(n4588), .CP(clock), .Q(result[23]) );
  CFD1QXL \result_reg[21]  ( .D(n4590), .CP(clock), .Q(result[21]) );
  CFD1QXL \result_reg[19]  ( .D(n4592), .CP(clock), .Q(result[19]) );
  CFD1QXL \result_reg[17]  ( .D(n4594), .CP(clock), .Q(result[17]) );
  CFD1QXL \result_reg[15]  ( .D(n4596), .CP(clock), .Q(result[15]) );
  CFD1QXL \result_reg[13]  ( .D(n4598), .CP(clock), .Q(result[13]) );
  CFD1QXL \result_reg[11]  ( .D(n4600), .CP(clock), .Q(result[11]) );
  CFD1QXL \result_reg[33]  ( .D(n4602), .CP(clock), .Q(result[33]) );
  CFD1QXL \result_reg[35]  ( .D(n4604), .CP(clock), .Q(result[35]) );
  CFD1QXL \result_reg[37]  ( .D(n4606), .CP(clock), .Q(result[37]) );
  CFD1QXL \result_reg[39]  ( .D(n4608), .CP(clock), .Q(result[39]) );
  CFD1QXL \result_reg[41]  ( .D(n4610), .CP(clock), .Q(result[41]) );
  CFD1QXL \result_reg[43]  ( .D(n4612), .CP(clock), .Q(result[43]) );
  CFD1QXL \result_reg[45]  ( .D(n4614), .CP(clock), .Q(result[45]) );
  CFD1QXL \result_reg[47]  ( .D(n4616), .CP(clock), .Q(result[47]) );
  CFD1QXL \result_reg[49]  ( .D(n4618), .CP(clock), .Q(result[49]) );
  CFD1QXL \result_reg[51]  ( .D(n4620), .CP(clock), .Q(result[51]) );
  CFD1QXL \result_reg[53]  ( .D(n4622), .CP(clock), .Q(result[53]) );
  CFD1QXL \result_reg[55]  ( .D(n4624), .CP(clock), .Q(result[55]) );
  CFD1QXL \result_reg[57]  ( .D(n4626), .CP(clock), .Q(result[57]) );
  CFD1QXL \result_reg[59]  ( .D(n4628), .CP(clock), .Q(result[59]) );
  CFD1QXL \result_reg[61]  ( .D(n4630), .CP(clock), .Q(result[61]) );
  CFD1QXL \result_reg[30]  ( .D(n4632), .CP(clock), .Q(result[30]) );
  CFD1QXL \result_reg[28]  ( .D(n4634), .CP(clock), .Q(result[28]) );
  CFD1QXL \result_reg[26]  ( .D(n4636), .CP(clock), .Q(result[26]) );
  CFD1QXL \result_reg[24]  ( .D(n4638), .CP(clock), .Q(result[24]) );
  CFD1QXL \result_reg[22]  ( .D(n4640), .CP(clock), .Q(result[22]) );
  CFD1QXL \result_reg[20]  ( .D(n4642), .CP(clock), .Q(result[20]) );
  CFD1QXL \result_reg[18]  ( .D(n4644), .CP(clock), .Q(result[18]) );
  CFD1QXL \result_reg[16]  ( .D(n4646), .CP(clock), .Q(result[16]) );
  CFD1QXL \result_reg[14]  ( .D(n4648), .CP(clock), .Q(result[14]) );
  CFD1QXL \result_reg[12]  ( .D(n4650), .CP(clock), .Q(result[12]) );
  CFD1QXL \result_reg[10]  ( .D(n4652), .CP(clock), .Q(result[10]) );
  CFD1QXL \result_reg[32]  ( .D(n4654), .CP(clock), .Q(result[32]) );
  CFD1QXL \result_reg[34]  ( .D(n4656), .CP(clock), .Q(result[34]) );
  CFD1QXL \result_reg[36]  ( .D(n4658), .CP(clock), .Q(result[36]) );
  CFD1QXL \result_reg[38]  ( .D(n4660), .CP(clock), .Q(result[38]) );
  CFD1QXL \result_reg[40]  ( .D(n4662), .CP(clock), .Q(result[40]) );
  CFD1QXL \result_reg[42]  ( .D(n4664), .CP(clock), .Q(result[42]) );
  CFD1QXL \result_reg[44]  ( .D(n4666), .CP(clock), .Q(result[44]) );
  CFD1QXL \result_reg[46]  ( .D(n4668), .CP(clock), .Q(result[46]) );
  CFD1QXL \result_reg[48]  ( .D(n4670), .CP(clock), .Q(result[48]) );
  CFD1QXL \result_reg[50]  ( .D(n4672), .CP(clock), .Q(result[50]) );
  CFD1QXL \result_reg[52]  ( .D(n4674), .CP(clock), .Q(result[52]) );
  CFD1QXL \result_reg[54]  ( .D(n4676), .CP(clock), .Q(result[54]) );
  CFD1QXL \result_reg[56]  ( .D(n4678), .CP(clock), .Q(result[56]) );
  CFD1QXL \result_reg[58]  ( .D(n4680), .CP(clock), .Q(result[58]) );
  CFD1QXL \result_reg[60]  ( .D(n4682), .CP(clock), .Q(result[60]) );
  CFD1QXL \result_reg[62]  ( .D(n4684), .CP(clock), .Q(result[62]) );
  CFD1QXL \result_copy_reg[60]  ( .D(n4686), .CP(clock), .Q(D[28]) );
  CFD1QXL \opera1_copy_reg[29]  ( .D(n4688), .CP(clock), .Q(opera1_copy[29])
         );
  CFD1QXL \opera1_copydiv_reg[31]  ( .D(n3105), .CP(clock), .Q(
        opera1_copydiv[31]) );
  CFD1QXL \result_copy_reg[62]  ( .D(n4691), .CP(clock), .Q(D[30]) );
  CFD1XL \opera1_copydiv_reg[29]  ( .D(n4693), .CP(clock), .QN(n1772) );
  CFD1XL \opera1_copydiv_reg[27]  ( .D(n4699), .CP(clock), .QN(
        \intadd_0/B[26] ) );
  CFD1QXL \result_not_reg[60]  ( .D(n4704), .CP(clock), .Q(result_not[60]) );
  CFD1QXL \result_not_reg[54]  ( .D(n4705), .CP(clock), .Q(result_not[54]) );
  CFD1QXL \result_not_reg[56]  ( .D(n4706), .CP(clock), .Q(result_not[56]) );
  CFD1QXL \result_not_reg[58]  ( .D(n4707), .CP(clock), .Q(result_not[58]) );
  CFD1XL \result_copy_reg[0]  ( .D(n1620), .CP(clock), .Q(n4488), .QN(n335) );
  CFD1QXL \result_copy_reg[63]  ( .D(n4709), .CP(clock), .Q(D[31]) );
  CFD1XL OPE_reg ( .D(n1622), .CP(clock), .Q(n4489), .QN(n1770) );
  CFD1QXL \opera1_copy_reg[25]  ( .D(n4711), .CP(clock), .Q(opera1_copy[25])
         );
  CFD1QXL \i_reg[27]  ( .D(n4714), .CP(clock), .Q(i[27]) );
  CFD1QXL \opera1_copy_reg[22]  ( .D(n4716), .CP(clock), .Q(opera1_copy[22])
         );
  CFD1QXL \opera1_copydiv_reg[20]  ( .D(n4718), .CP(clock), .Q(
        opera1_copydiv[20]) );
  CFD1QXL \opera1_copydiv_reg[22]  ( .D(n4722), .CP(clock), .Q(
        opera1_copydiv[22]) );
  CFD1QXL \opera1_copydiv_reg[24]  ( .D(n4724), .CP(clock), .Q(
        opera1_copydiv[24]) );
  CFD1QXL \opera1_copy_reg[21]  ( .D(n4726), .CP(clock), .Q(opera1_copy[21])
         );
  CFD1QXL \opera1_copy_reg[24]  ( .D(n4727), .CP(clock), .Q(opera1_copy[24])
         );
  CFD1QXL \opera1_copy_reg[23]  ( .D(n4732), .CP(clock), .Q(opera1_copy[23])
         );
  CFD1QXL \opera1_copy_reg[20]  ( .D(n4735), .CP(clock), .Q(opera1_copy[20])
         );
  CFD1QXL \opera1_copy_reg[19]  ( .D(n4739), .CP(clock), .Q(opera1_copy[19])
         );
  CFD1QXL \i_reg[30]  ( .D(n4741), .CP(clock), .Q(i[30]) );
  CFD1QXL \i_reg[22]  ( .D(n4743), .CP(clock), .Q(i[22]) );
  CFD1QXL \i_reg[14]  ( .D(n4745), .CP(clock), .Q(i[14]) );
  CFD1QXL \i_reg[8]  ( .D(n4747), .CP(clock), .Q(i[8]) );
  CFD1QXL \i_reg[6]  ( .D(n4749), .CP(clock), .Q(i[6]) );
  CFD1QXL \i_reg[16]  ( .D(n4751), .CP(clock), .Q(i[16]) );
  CFD1QXL \i_reg[18]  ( .D(n4753), .CP(clock), .Q(i[18]) );
  CFD1QXL \i_reg[20]  ( .D(n4755), .CP(clock), .Q(i[20]) );
  CFD1QXL \i_reg[28]  ( .D(n4757), .CP(clock), .Q(i[28]) );
  CFD1QXL \i_reg[24]  ( .D(n4759), .CP(clock), .Q(i[24]) );
  CFD1QXL \i_reg[26]  ( .D(n4761), .CP(clock), .Q(i[26]) );
  CFD1QXL \i_reg[10]  ( .D(n4763), .CP(clock), .Q(i[10]) );
  CFD1QXL \i_reg[12]  ( .D(n4765), .CP(clock), .Q(i[12]) );
  CFD1QXL \i_reg[29]  ( .D(n4767), .CP(clock), .Q(i[29]) );
  CFD1QXL \i_reg[7]  ( .D(n4769), .CP(clock), .Q(i[7]) );
  CFD1QXL \i_reg[17]  ( .D(n4771), .CP(clock), .Q(i[17]) );
  CFD1QXL \i_reg[9]  ( .D(n4773), .CP(clock), .Q(i[9]) );
  CFD1QXL \i_reg[25]  ( .D(n4775), .CP(clock), .Q(i[25]) );
  CFD1QXL \i_reg[13]  ( .D(n4777), .CP(clock), .Q(i[13]) );
  CFD1QXL \i_reg[23]  ( .D(n4779), .CP(clock), .Q(i[23]) );
  CFD1QXL \i_reg[11]  ( .D(n4781), .CP(clock), .Q(i[11]) );
  CFD1QXL \i_reg[15]  ( .D(n4783), .CP(clock), .Q(i[15]) );
  CFD1QXL \i_reg[21]  ( .D(n4785), .CP(clock), .Q(i[21]) );
  CFD1QXL \i_reg[19]  ( .D(n4787), .CP(clock), .Q(i[19]) );
  CFD1QXL \i_reg[1]  ( .D(n4789), .CP(clock), .Q(i[1]) );
  CFD1QXL \i_reg[2]  ( .D(n4790), .CP(clock), .Q(i[2]) );
  CFD1QXL \i_reg[0]  ( .D(n4792), .CP(clock), .Q(i[0]) );
  CFD1QXL \result_copy_reg[56]  ( .D(n4795), .CP(clock), .Q(D[24]) );
  CFD1QXL \result_copy_reg[52]  ( .D(n4797), .CP(clock), .Q(D[20]) );
  CFD1QXL \i_reg[5]  ( .D(n1623), .CP(clock), .Q(i[5]) );
  CFD1QXL \i_reg[3]  ( .D(n4799), .CP(clock), .Q(i[3]) );
  CFD1QXL \result_copy_reg[58]  ( .D(n4801), .CP(clock), .Q(D[26]) );
  CFD1QXL \result_copy_reg[54]  ( .D(n4805), .CP(clock), .Q(D[22]) );
  CFD1QXL \i_reg[4]  ( .D(n4809), .CP(clock), .Q(i[4]) );
  CFD1XL \opera1_copydiv_reg[25]  ( .D(n4810), .CP(clock), .QN(
        \intadd_0/B[24] ) );
  CFD1XL \opera1_copydiv_reg[21]  ( .D(n4813), .CP(clock), .QN(
        \intadd_0/B[20] ) );
  CFD1XL \opera1_copydiv_reg[23]  ( .D(n4819), .CP(clock), .QN(
        \intadd_0/B[22] ) );
  CFD1QXL \result_not_reg[46]  ( .D(n4822), .CP(clock), .Q(result_not[46]) );
  CFD1QXL \result_not_reg[48]  ( .D(n4823), .CP(clock), .Q(result_not[48]) );
  CFD1QXL \result_not_reg[50]  ( .D(n4824), .CP(clock), .Q(result_not[50]) );
  CFD1QXL \result_not_reg[52]  ( .D(n4825), .CP(clock), .Q(result_not[52]) );
  CFD1QXL \result_not_reg[44]  ( .D(n4826), .CP(clock), .Q(result_not[44]) );
  CFD2QXL \cust_reg[1]  ( .D(N145), .CP(clock), .CD(n3076), .Q(\cust[1] ) );
  CFD1QXL \opera1_copy_reg[18]  ( .D(n4830), .CP(clock), .Q(opera1_copy[18])
         );
  CFD1QXL \opera1_copy_reg[14]  ( .D(n4833), .CP(clock), .Q(opera1_copy[14])
         );
  CFD1QXL \opera1_copydiv_reg[14]  ( .D(n4838), .CP(clock), .Q(
        opera1_copydiv[14]) );
  CFD1QXL \opera1_copydiv_reg[16]  ( .D(n4839), .CP(clock), .Q(
        opera1_copydiv[16]) );
  CFD1QXL \opera1_copydiv_reg[18]  ( .D(n4843), .CP(clock), .Q(
        opera1_copydiv[18]) );
  CFD1QXL \opera1_copy_reg[17]  ( .D(n4844), .CP(clock), .Q(opera1_copy[17])
         );
  CFD1QXL \opera1_copy_reg[13]  ( .D(n4846), .CP(clock), .Q(opera1_copy[13])
         );
  CFD1QXL \opera1_copy_reg[16]  ( .D(n4848), .CP(clock), .Q(opera1_copy[16])
         );
  CFD1QXL \opera1_copy_reg[15]  ( .D(n4849), .CP(clock), .Q(opera1_copy[15])
         );
  CFD1QXL \result_copy_reg[48]  ( .D(n4850), .CP(clock), .Q(D[16]) );
  CFD1QXL \result_copy_reg[50]  ( .D(n4852), .CP(clock), .Q(D[18]) );
  CFD1QXL \result_copy_reg[46]  ( .D(n4856), .CP(clock), .Q(D[14]) );
  CFD1XL \opera1_copydiv_reg[13]  ( .D(n4860), .CP(clock), .QN(
        \intadd_0/B[12] ) );
  CFD1XL \opera1_copydiv_reg[17]  ( .D(n4864), .CP(clock), .QN(
        \intadd_0/B[16] ) );
  CFD1XL \opera1_copydiv_reg[19]  ( .D(n4869), .CP(clock), .QN(
        \intadd_0/B[18] ) );
  CFD1XL \opera1_copydiv_reg[15]  ( .D(n4874), .CP(clock), .QN(
        \intadd_0/B[14] ) );
  CFD1QXL \result_not_reg[36]  ( .D(n4880), .CP(clock), .Q(result_not[36]) );
  CFD1QXL \result_not_reg[38]  ( .D(n4881), .CP(clock), .Q(result_not[38]) );
  CFD1QXL \result_not_reg[40]  ( .D(n4882), .CP(clock), .Q(result_not[40]) );
  CFD1QXL \result_not_reg[42]  ( .D(n4883), .CP(clock), .Q(result_not[42]) );
  CFD1QXL \opera1_copy_reg[12]  ( .D(n4884), .CP(clock), .Q(opera1_copy[12])
         );
  CFD1QXL \opera1_copy_reg[10]  ( .D(n4887), .CP(clock), .Q(opera1_copy[10])
         );
  CFD1QXL \opera1_copy_reg[6]  ( .D(n4890), .CP(clock), .Q(opera1_copy[6]) );
  CFD1QXL \opera1_copydiv_reg[8]  ( .D(n4893), .CP(clock), .Q(
        opera1_copydiv[8]) );
  CFD1QXL \opera1_copydiv_reg[10]  ( .D(n4897), .CP(clock), .Q(
        opera1_copydiv[10]) );
  CFD1QXL \opera1_copydiv_reg[12]  ( .D(n4898), .CP(clock), .Q(
        opera1_copydiv[12]) );
  CFD1QXL \opera1_copy_reg[9]  ( .D(n4903), .CP(clock), .Q(opera1_copy[9]) );
  CFD1QXL \opera1_copy_reg[11]  ( .D(n4905), .CP(clock), .Q(opera1_copy[11])
         );
  CFD1QXL \opera1_copy_reg[8]  ( .D(n4907), .CP(clock), .Q(opera1_copy[8]) );
  CFD1QXL \opera1_copy_reg[7]  ( .D(n4908), .CP(clock), .Q(opera1_copy[7]) );
  CFD1QXL \result_copy_reg[44]  ( .D(n4909), .CP(clock), .Q(D[12]) );
  CFD1QXL \result_copy_reg[40]  ( .D(n4911), .CP(clock), .Q(D[8]) );
  CFD1QXL \result_copy_reg[42]  ( .D(n4913), .CP(clock), .Q(D[10]) );
  CFD1XL \opera1_copydiv_reg[9]  ( .D(n4917), .CP(clock), .QN(\intadd_0/B[8] )
         );
  CFD1XL \opera1_copydiv_reg[7]  ( .D(n4922), .CP(clock), .QN(\intadd_0/B[6] )
         );
  CFD1XL \opera1_copydiv_reg[11]  ( .D(n4927), .CP(clock), .QN(
        \intadd_0/B[10] ) );
  CFD1QXL \result_not_reg[34]  ( .D(n4932), .CP(clock), .Q(result_not[34]) );
  CFD1QXL \result_not_reg[30]  ( .D(n4933), .CP(clock), .Q(result_not[30]) );
  CFD1QXL \result_not_reg[32]  ( .D(n1522), .CP(clock), .Q(result_not[32]) );
  CFD1QXL \result_not_reg[28]  ( .D(n4934), .CP(clock), .Q(result_not[28]) );
  CFD1QXL \opera1_copydiv_reg[6]  ( .D(n4937), .CP(clock), .Q(
        opera1_copydiv[6]) );
  CFD1QXL \opera1_copy_reg[2]  ( .D(n4939), .CP(clock), .Q(opera1_copy[2]) );
  CFD1QXL \opera1_copydiv_reg[2]  ( .D(n4942), .CP(clock), .Q(
        opera1_copydiv[2]) );
  CFD1QXL \opera1_copydiv_reg[4]  ( .D(n4947), .CP(clock), .Q(
        opera1_copydiv[4]) );
  CFD1QXL \opera1_copy_reg[5]  ( .D(n4949), .CP(clock), .Q(opera1_copy[5]) );
  CFD1QXL \opera1_copy_reg[4]  ( .D(n4951), .CP(clock), .Q(opera1_copy[4]) );
  CFD1QXL \opera1_copy_reg[3]  ( .D(n4954), .CP(clock), .Q(opera1_copy[3]) );
  CFD1QXL \opera1_copy_reg[1]  ( .D(n4955), .CP(clock), .Q(opera1_copy[1]) );
  CFD1QXL \opera1_copydiv_reg[0]  ( .D(n4956), .CP(clock), .Q(
        opera1_copydiv[0]) );
  CFD1QXL \result_copy_reg[34]  ( .D(n4957), .CP(clock), .Q(D[2]) );
  CFD1QXL \result_copy_reg[38]  ( .D(n4961), .CP(clock), .Q(D[6]) );
  CFD1XL \opera1_copydiv_reg[5]  ( .D(n4965), .CP(clock), .QN(\intadd_0/B[4] )
         );
  CFD1XL \opera1_copydiv_reg[1]  ( .D(n4970), .CP(clock), .QN(\intadd_0/B[0] )
         );
  CFD1XL \opera1_copydiv_reg[3]  ( .D(n4975), .CP(clock), .QN(\intadd_0/B[2] )
         );
  CFD1QXL \result_not_reg[26]  ( .D(n4978), .CP(clock), .Q(result_not[26]) );
  CFD1QXL \result_not_reg[24]  ( .D(n4979), .CP(clock), .Q(result_not[24]) );
  CFD1QXL \result_not_reg[22]  ( .D(n4980), .CP(clock), .Q(result_not[22]) );
  CFD1QXL \result_not_reg[20]  ( .D(n4981), .CP(clock), .Q(result_not[20]) );
  CFD1QXL \result_not_reg[18]  ( .D(n4982), .CP(clock), .Q(result_not[18]) );
  CFD1QXL \opera1_copy_reg[0]  ( .D(n4983), .CP(clock), .Q(opera1_copy[0]) );
  CFD1QXL \result_copy_reg[32]  ( .D(n4989), .CP(clock), .Q(D[0]) );
  CFD1XL \result_copy_reg[36]  ( .D(n4993), .CP(clock), .QN(n1741) );
  CFD1QXL \result_not_reg[16]  ( .D(n4995), .CP(clock), .Q(result_not[16]) );
  CFD1QXL \result_not_reg[14]  ( .D(n4996), .CP(clock), .Q(result_not[14]) );
  CFD1QXL \result_not_reg[12]  ( .D(n4997), .CP(clock), .Q(result_not[12]) );
  CFD1QXL \result_not_reg[10]  ( .D(n4998), .CP(clock), .Q(result_not[10]) );
  CFD1QXL w4_reg ( .D(n4999), .CP(clock), .Q(w4) );
  CFD1QXL \result_not_reg[8]  ( .D(n5000), .CP(clock), .Q(result_not[8]) );
  CFD1QXL \result_not_reg[4]  ( .D(n5001), .CP(clock), .Q(result_not[4]) );
  CFD1QXL \result_not_reg[0]  ( .D(n1554), .CP(clock), .Q(result_not[0]) );
  CFD1QXL \result_not_reg[6]  ( .D(n5002), .CP(clock), .Q(result_not[6]) );
  CFD1QXL \result_not_reg[2]  ( .D(n5003), .CP(clock), .Q(result_not[2]) );
  CFD4XL \cust_reg[2]  ( .D(n5004), .CP(clock), .SD(n3076), .Q(n284), .QN(
        n3479) );
  CFD4XL \cust_reg[0]  ( .D(n259), .CP(clock), .SD(n3076), .Q(n260), .QN(n4472) );
  CFD1QXL \result_not_reg[31]  ( .D(n5011), .CP(clock), .Q(result_not[31]) );
  CFD1QXL \result_not_reg[29]  ( .D(n5012), .CP(clock), .Q(result_not[29]) );
  CFD1QXL \result_not_reg[27]  ( .D(n5013), .CP(clock), .Q(result_not[27]) );
  CFD1QXL \result_not_reg[25]  ( .D(n5014), .CP(clock), .Q(result_not[25]) );
  CFD1QXL \result_not_reg[23]  ( .D(n5015), .CP(clock), .Q(result_not[23]) );
  CFD1QXL \result_not_reg[21]  ( .D(n5016), .CP(clock), .Q(result_not[21]) );
  CFD1QXL \result_not_reg[19]  ( .D(n5017), .CP(clock), .Q(result_not[19]) );
  CFD1QXL \result_not_reg[17]  ( .D(n5018), .CP(clock), .Q(result_not[17]) );
  CFD1QXL \result_not_reg[15]  ( .D(n5019), .CP(clock), .Q(result_not[15]) );
  CFD1QXL \result_not_reg[13]  ( .D(n5020), .CP(clock), .Q(result_not[13]) );
  CFD1QXL \result_not_reg[11]  ( .D(n5021), .CP(clock), .Q(result_not[11]) );
  CFD1QXL \result_not_reg[9]  ( .D(n5022), .CP(clock), .Q(result_not[9]) );
  CFD1QXL \result_not_reg[7]  ( .D(n5023), .CP(clock), .Q(result_not[7]) );
  CFD1QXL \result_not_reg[5]  ( .D(n5025), .CP(clock), .Q(result_not[5]) );
  CFD1QXL \result_not_reg[3]  ( .D(n5026), .CP(clock), .Q(result_not[3]) );
  CFD1QXL \result_not_reg[1]  ( .D(n5028), .CP(clock), .Q(result_not[1]) );
  CFD1QXL \result_not_reg[37]  ( .D(n5030), .CP(clock), .Q(result_not[37]) );
  CFD1QXL \result_not_reg[35]  ( .D(n5031), .CP(clock), .Q(result_not[35]) );
  CFD1QXL \result_not_reg[33]  ( .D(n5032), .CP(clock), .Q(result_not[33]) );
  CFD1QXL \result_not_reg[39]  ( .D(n5033), .CP(clock), .Q(result_not[39]) );
  CFD1QXL \result_copy_reg[9]  ( .D(n5034), .CP(clock), .Q(result_copy[9]) );
  CFD1QXL \result_copy_reg[5]  ( .D(n5037), .CP(clock), .Q(result_copy[5]) );
  CFD1QXL \result_copy_reg[1]  ( .D(n5042), .CP(clock), .Q(result_copy[1]) );
  CFD1QXL \result_not_reg[41]  ( .D(n5048), .CP(clock), .Q(result_not[41]) );
  CFD1QXL \result_copy_reg[13]  ( .D(n5049), .CP(clock), .Q(result_copy[13])
         );
  CFD1QXL \result_not_reg[43]  ( .D(n5054), .CP(clock), .Q(result_not[43]) );
  CFD1QXL \result_copy_reg[15]  ( .D(n5055), .CP(clock), .Q(n4469) );
  CFD1QXL \result_copy_reg[17]  ( .D(n5060), .CP(clock), .Q(result_copy[17])
         );
  CFD1QXL \result_copy_reg[19]  ( .D(n5065), .CP(clock), .Q(result_copy[19])
         );
  CFD1QXL \result_not_reg[45]  ( .D(n5070), .CP(clock), .Q(result_not[45]) );
  CFD1QXL \result_copy_reg[21]  ( .D(n5071), .CP(clock), .Q(result_copy[21])
         );
  CFD1QXL \result_copy_reg[23]  ( .D(n5076), .CP(clock), .Q(result_copy[23])
         );
  CFD1QXL \result_not_reg[47]  ( .D(n5081), .CP(clock), .Q(result_not[47]) );
  CFD1QXL \result_copy_reg[25]  ( .D(n5082), .CP(clock), .Q(result_copy[25])
         );
  CFD1QXL \result_copy_reg[27]  ( .D(n5087), .CP(clock), .Q(result_copy[27])
         );
  CFD1QXL \result_not_reg[49]  ( .D(n5092), .CP(clock), .Q(result_not[49]) );
  CFD1QXL \result_copy_reg[29]  ( .D(n5093), .CP(clock), .Q(result_copy[29])
         );
  CFD1QXL \result_not_reg[51]  ( .D(n5098), .CP(clock), .Q(result_not[51]) );
  CFD1QXL \result_copy_reg[31]  ( .D(n5099), .CP(clock), .Q(result_copy[31])
         );
  CFD1QXL \result_not_reg[53]  ( .D(n5103), .CP(clock), .Q(result_not[53]) );
  CFD1QXL \result_not_reg[55]  ( .D(n5104), .CP(clock), .Q(result_not[55]) );
  CFD1QXL \result_not_reg[57]  ( .D(n5105), .CP(clock), .Q(result_not[57]) );
  CFD1QXL \result_not_reg[59]  ( .D(n5106), .CP(clock), .Q(result_not[59]) );
  CFD1QXL \result_not_reg[61]  ( .D(n5107), .CP(clock), .Q(result_not[61]) );
  CFD1XL valid_reg ( .D(n5108), .CP(clock), .Q(valid), .QN(n3389) );
  CFD1XL \result_copy_reg[33]  ( .D(n5109), .CP(clock), .Q(n1773), .QN(n3316)
         );
  CFD1XL \result_copy_reg[35]  ( .D(n5114), .CP(clock), .Q(n1796), .QN(n3272)
         );
  CFD1XL \result_copy_reg[37]  ( .D(n5115), .CP(clock), .Q(n1797), .QN(n3266)
         );
  CFD1XL \result_copy_reg[39]  ( .D(n5118), .CP(clock), .Q(n1798), .QN(n3261)
         );
  CFD1XL \result_copy_reg[41]  ( .D(n5121), .CP(clock), .Q(n1799), .QN(n3256)
         );
  CFD1XL \result_copy_reg[43]  ( .D(n5124), .CP(clock), .Q(n1800), .QN(n3251)
         );
  CFD1XL \result_copy_reg[45]  ( .D(n5128), .CP(clock), .Q(n1801), .QN(n3246)
         );
  CFD1XL \result_copy_reg[47]  ( .D(n5131), .CP(clock), .Q(n1802), .QN(n3241)
         );
  CFD1XL \result_copy_reg[49]  ( .D(n5134), .CP(clock), .Q(n1803), .QN(n3236)
         );
  CFD1XL \result_copy_reg[51]  ( .D(n5137), .CP(clock), .Q(n1804), .QN(n3231)
         );
  CFD1XL \result_copy_reg[53]  ( .D(n5140), .CP(clock), .Q(n1805), .QN(n3226)
         );
  CFD1XL \result_copy_reg[55]  ( .D(n5143), .CP(clock), .Q(n1806), .QN(n3221)
         );
  CFD1XL \result_copy_reg[57]  ( .D(n5147), .CP(clock), .Q(n1807), .QN(n3216)
         );
  CFD1XL \result_copy_reg[59]  ( .D(n5150), .CP(clock), .Q(n1808), .QN(n3211)
         );
  CFD1XL \result_copy_reg[61]  ( .D(n5154), .CP(clock), .Q(n1734), .QN(n3397)
         );
  COND3X2 U3289 ( .A(n327), .B(n3772), .C(n3824), .D(n3825), .Z(n1610) );
  CNIVXL U3290 ( .A(opera2[0]), .Z(n4708) );
  CNIVX1 U3291 ( .A(n3198), .Z(n4470) );
  CNIVX1 U3292 ( .A(n4473), .Z(n4471) );
  CNR3X1 U3293 ( .A(n3758), .B(n3944), .C(n4489), .Z(n5179) );
  CNR3X1 U3294 ( .A(n3944), .B(n1770), .C(n3758), .Z(n5178) );
  CND2X1 U3295 ( .A(n4472), .B(n3414), .Z(n3758) );
  CNR2X1 U3296 ( .A(n4472), .B(\cust[1] ), .Z(n3751) );
  CANR11X1 U3297 ( .A(n4470), .B(n3774), .C(n3777), .D(n3757), .Z(n3769) );
  CAN3X2 U3298 ( .A(n3768), .B(n3769), .C(n3770), .Z(n4473) );
  CIVX2 U3299 ( .A(n4471), .Z(n1620) );
  CIVDXL U3300 ( .A(n4309), .Z0(n4474), .Z1(n4475) );
  CIVDX1 U3301 ( .A(n3483), .Z0(n4476), .Z1(n4477) );
  CIVDX1 U3302 ( .A(opera2[63]), .Z0(n4478), .Z1(n4479) );
  CIVDX1 U3303 ( .A(n3647), .Z0(n4480), .Z1(n4481) );
  CIVDXL U3304 ( .A(n3753), .Z0(n4482), .Z1(n4483) );
  CIVX2 U3305 ( .A(n4486), .Z(n5192) );
  CAN2X1 U3306 ( .A(n4179), .B(n1770), .Z(n4484) );
  CIVXL U3307 ( .A(n327), .Z(n3377) );
  CANR2X2 U3308 ( .A(result_not[5]), .B(n4168), .C(n332), .D(n4179), .Z(n4183)
         );
  CANR2X2 U3309 ( .A(result_not[9]), .B(n4168), .C(n329), .D(n4179), .Z(n4187)
         );
  COR2X1 U3310 ( .A(n4488), .B(n3772), .Z(n4485) );
  COR2X1 U3311 ( .A(n4476), .B(n3136), .Z(n4486) );
  CIVX2 U3312 ( .A(n5157), .Z(n5189) );
  COR2X1 U3313 ( .A(n3772), .B(n335), .Z(n4487) );
  CND4XL U3314 ( .A(n4137), .B(n4138), .C(n4139), .D(n5155), .Z(n1559) );
  CND2XL U3315 ( .A(n3751), .B(n3479), .Z(n4170) );
  CNIVXL U3316 ( .A(reset), .Z(n4794) );
  CAN4XL U3317 ( .A(n4476), .B(n5186), .C(n3754), .D(n4172), .Z(n3648) );
  COND3XL U3318 ( .A(n3201), .B(n4143), .C(n4272), .D(n4273), .Z(n1491) );
  CNIVX1 U3319 ( .A(n1491), .Z(n4490) );
  CNIVXL U3320 ( .A(opera2[3]), .Z(n4494) );
  CNIVX1 U3321 ( .A(n4494), .Z(n4491) );
  CNIVX1 U3322 ( .A(n4493), .Z(n4492) );
  CNIVX1 U3323 ( .A(n4495), .Z(n4493) );
  CNIVX1 U3324 ( .A(n1617), .Z(n4495) );
  CANR2XL U3325 ( .A(n5182), .B(n3794), .C(n5180), .D(n4491), .Z(n3792) );
  CNIVXL U3326 ( .A(opera2[7]), .Z(n4499) );
  CNIVX1 U3327 ( .A(n4499), .Z(n4496) );
  CNIVX1 U3328 ( .A(n4498), .Z(n4497) );
  CNIVX1 U3329 ( .A(n4500), .Z(n4498) );
  CNIVX1 U3330 ( .A(n1613), .Z(n4500) );
  CANR2XL U3331 ( .A(n5182), .B(n3813), .C(n5180), .D(n4496), .Z(n3811) );
  CDLY1XL U3332 ( .A(n1594), .Z(n4502) );
  CNIVX1 U3333 ( .A(opera2[26]), .Z(n4501) );
  CANR2XL U3334 ( .A(n3908), .B(n3909), .C(n5180), .D(n4501), .Z(n3906) );
  CDLY1XL U3335 ( .A(n1608), .Z(n4504) );
  COND3XL U3336 ( .A(n3772), .B(n3288), .C(n3833), .D(n3834), .Z(n1608) );
  CNIVX1 U3337 ( .A(opera2[12]), .Z(n4503) );
  CANR2XL U3338 ( .A(n3835), .B(n3836), .C(n5180), .D(n4503), .Z(n3833) );
  CDLY1XL U3339 ( .A(n1604), .Z(n4506) );
  COND3XL U3340 ( .A(n3772), .B(n3287), .C(n3854), .D(n3855), .Z(n1604) );
  CNIVX1 U3341 ( .A(opera2[16]), .Z(n4505) );
  CANR2XL U3342 ( .A(n3856), .B(n3857), .C(n5180), .D(n4505), .Z(n3854) );
  CDLY1XL U3343 ( .A(n1596), .Z(n4508) );
  COND3XL U3344 ( .A(n3772), .B(n3286), .C(n3896), .D(n3897), .Z(n1596) );
  CNIVX1 U3345 ( .A(opera2[24]), .Z(n4507) );
  CANR2XL U3346 ( .A(n3898), .B(n3899), .C(n5180), .D(n4507), .Z(n3896) );
  CDLY1XL U3347 ( .A(opera2[10]), .Z(n4509) );
  CNIVX1 U3348 ( .A(n1610), .Z(n4510) );
  CANR2XL U3349 ( .A(n3826), .B(n3778), .C(n5180), .D(n4509), .Z(n3824) );
  CDLY1XL U3350 ( .A(n1606), .Z(n4512) );
  CNIVX1 U3351 ( .A(opera2[14]), .Z(n4511) );
  CANR2XL U3352 ( .A(n3845), .B(n3846), .C(n5180), .D(n4511), .Z(n3843) );
  CDLY1XL U3353 ( .A(n1602), .Z(n4514) );
  CNIVX1 U3354 ( .A(opera2[18]), .Z(n4513) );
  CANR2XL U3355 ( .A(n3866), .B(n3867), .C(n5180), .D(n4513), .Z(n3864) );
  CDLY1XL U3356 ( .A(n1600), .Z(n4516) );
  COND3XL U3357 ( .A(n3772), .B(n3294), .C(n3875), .D(n3876), .Z(n1600) );
  CNIVX1 U3358 ( .A(opera2[20]), .Z(n4515) );
  CANR2XL U3359 ( .A(n3877), .B(n3878), .C(n5180), .D(n4515), .Z(n3875) );
  CDLY1XL U3360 ( .A(n1598), .Z(n4518) );
  CNIVX1 U3361 ( .A(opera2[22]), .Z(n4517) );
  CANR2XL U3362 ( .A(n3887), .B(n3888), .C(n5180), .D(n4517), .Z(n3885) );
  CDLY1XL U3363 ( .A(n1592), .Z(n4520) );
  COND3XL U3364 ( .A(n3772), .B(n3293), .C(n3917), .D(n3918), .Z(n1592) );
  CNIVX1 U3365 ( .A(opera2[28]), .Z(n4519) );
  CANR2XL U3366 ( .A(n3919), .B(n3920), .C(n5180), .D(n4519), .Z(n3917) );
  CDLY1XL U3367 ( .A(n1614), .Z(n4522) );
  COND3XL U3368 ( .A(n3772), .B(n3365), .C(n3805), .D(n3806), .Z(n1614) );
  CNIVX1 U3369 ( .A(opera2[6]), .Z(n4521) );
  CANR2XL U3370 ( .A(n3807), .B(n3808), .C(n5180), .D(n4521), .Z(n3805) );
  CND2XL U3371 ( .A(n3786), .B(n4162), .Z(n3790) );
  CNIVXL U3372 ( .A(opera2[2]), .Z(n4526) );
  CNIVX1 U3373 ( .A(n4525), .Z(n4523) );
  CNIVX1 U3374 ( .A(n4526), .Z(n4524) );
  CNIVX1 U3375 ( .A(n1618), .Z(n4525) );
  CANR2XL U3376 ( .A(n3789), .B(n3790), .C(n5180), .D(n4524), .Z(n3787) );
  CNIVX1 U3377 ( .A(n1492), .Z(n4527) );
  CDLY1XL U3378 ( .A(n1590), .Z(n4529) );
  CNIVX1 U3379 ( .A(opera2[30]), .Z(n4528) );
  CANR2XL U3380 ( .A(n3929), .B(n3930), .C(n5180), .D(n4528), .Z(n3927) );
  CNIVXL U3381 ( .A(opera2[4]), .Z(n4533) );
  CNIVX1 U3382 ( .A(n4533), .Z(n4530) );
  CNIVX1 U3383 ( .A(n4532), .Z(n4531) );
  CNIVX1 U3384 ( .A(n4534), .Z(n4532) );
  CNIVX1 U3385 ( .A(n1616), .Z(n4534) );
  CANR2XL U3386 ( .A(n3798), .B(n5181), .C(n5180), .D(n4530), .Z(n3796) );
  COND3XL U3387 ( .A(n3772), .B(n3289), .C(n4536), .D(n3816), .Z(n1612) );
  CNIVX1 U3388 ( .A(n4538), .Z(n4535) );
  CNIVX1 U3389 ( .A(n4537), .Z(n4536) );
  CNIVX1 U3390 ( .A(n3815), .Z(n4537) );
  CNIVX1 U3391 ( .A(n1612), .Z(n4538) );
  CDLY1XL U3392 ( .A(n1609), .Z(n4540) );
  COND3XL U3393 ( .A(n3772), .B(n3367), .C(n3829), .D(n3830), .Z(n1609) );
  CNIVX1 U3394 ( .A(opera2[11]), .Z(n4539) );
  CANR2XL U3395 ( .A(n5182), .B(n3831), .C(n5180), .D(n4539), .Z(n3829) );
  CAOR1X4 U3396 ( .A(n4542), .B(n3078), .C(n4303), .Z(n1481) );
  CNIVX1 U3397 ( .A(n1481), .Z(n4541) );
  CNIVX1 U3398 ( .A(result[9]), .Z(n4542) );
  CAOR1X4 U3399 ( .A(n4544), .B(n3078), .C(n4298), .Z(n1483) );
  CNIVX1 U3400 ( .A(n1483), .Z(n4543) );
  CNIVX1 U3401 ( .A(result[7]), .Z(n4544) );
  CAOR1X4 U3402 ( .A(n4546), .B(n3078), .C(n4293), .Z(n1485) );
  CNIVX1 U3403 ( .A(n1485), .Z(n4545) );
  CNIVX1 U3404 ( .A(result[5]), .Z(n4546) );
  CAOR1X4 U3405 ( .A(n4548), .B(n3078), .C(n4288), .Z(n1487) );
  CNIVX1 U3406 ( .A(n1487), .Z(n4547) );
  CNIVX1 U3407 ( .A(result[3]), .Z(n4548) );
  CAOR1X4 U3408 ( .A(n4550), .B(n3078), .C(n4283), .Z(n1489) );
  CNIVX1 U3409 ( .A(n1489), .Z(n4549) );
  CNIVX1 U3410 ( .A(result[1]), .Z(n4550) );
  CAOR1X4 U3411 ( .A(n4552), .B(n3078), .C(n4296), .Z(n1484) );
  CNIVX1 U3412 ( .A(n1484), .Z(n4551) );
  CNIVX1 U3413 ( .A(result[6]), .Z(n4552) );
  CAOR1X4 U3414 ( .A(n4554), .B(n3078), .C(n4286), .Z(n1488) );
  CNIVX1 U3415 ( .A(n1488), .Z(n4553) );
  CNIVX1 U3416 ( .A(result[2]), .Z(n4554) );
  CAOR1X4 U3417 ( .A(n4556), .B(n3078), .C(n4280), .Z(n1490) );
  CNIVX1 U3418 ( .A(n1490), .Z(n4555) );
  CNIVX1 U3419 ( .A(result[0]), .Z(n4556) );
  CAOR1X4 U3420 ( .A(n4558), .B(n3078), .C(n4466), .Z(n1427) );
  CNIVX1 U3421 ( .A(n1427), .Z(n4557) );
  CNIVX1 U3422 ( .A(result[63]), .Z(n4558) );
  CAOR1X4 U3423 ( .A(n4560), .B(n3078), .C(n4301), .Z(n1482) );
  CNIVX1 U3424 ( .A(n1482), .Z(n4559) );
  CNIVX1 U3425 ( .A(result[8]), .Z(n4560) );
  CAOR1X4 U3426 ( .A(n4562), .B(n3078), .C(n4291), .Z(n1486) );
  CNIVX1 U3427 ( .A(n1486), .Z(n4561) );
  CNIVX1 U3428 ( .A(result[4]), .Z(n4562) );
  COND3XL U3429 ( .A(n3380), .B(n4477), .C(n3490), .D(n3491), .Z(n255) );
  CNIVX1 U3430 ( .A(n255), .Z(n4563) );
  COND4CXL U3431 ( .A(n3492), .B(n3489), .C(n3493), .D(n3137), .Z(n3491) );
  COND4CXL U3432 ( .A(n3487), .B(n4477), .C(n3494), .D(n4690), .Z(n3490) );
  CIVXL U3433 ( .A(muordi), .Z(n3200) );
  COND3XL U3434 ( .A(n3381), .B(n4477), .C(n3498), .D(n3499), .Z(n253) );
  CNIVX1 U3435 ( .A(n4565), .Z(n4564) );
  CNIVX1 U3436 ( .A(n253), .Z(n4565) );
  CNIVX1 U3437 ( .A(n4567), .Z(n4566) );
  CNIVXL U3438 ( .A(opera1[25]), .Z(n4812) );
  CNIVX1 U3439 ( .A(n251), .Z(n4567) );
  COND3X2 U3440 ( .A(n3382), .B(n4477), .C(n3510), .D(n3511), .Z(n251) );
  CIVXL U3441 ( .A(opera1_copydiv[26]), .Z(n3383) );
  CNIVX1 U3442 ( .A(n4569), .Z(n4568) );
  CNIVX1 U3443 ( .A(n4702), .Z(n4569) );
  CNIVX1 U3444 ( .A(n1660), .Z(n4570) );
  CIVXL U3445 ( .A(opera1_copydiv[28]), .Z(n3384) );
  CNIVX1 U3446 ( .A(n4572), .Z(n4571) );
  CNIVX1 U3447 ( .A(n4697), .Z(n4572) );
  CNIVX1 U3448 ( .A(n1658), .Z(n4573) );
  CNIVX1 U3449 ( .A(n4575), .Z(n4574) );
  CNIVX1 U3450 ( .A(n1656), .Z(n4575) );
  COND3XL U3451 ( .A(n3388), .B(n4477), .C(n3506), .D(n3507), .Z(n252) );
  CNIVX1 U3452 ( .A(n4577), .Z(n4576) );
  CNIVX1 U3453 ( .A(n4578), .Z(n4577) );
  CNIVX1 U3454 ( .A(n252), .Z(n4578) );
  COND3XL U3455 ( .A(n4477), .B(n3390), .C(n3484), .D(n3485), .Z(n256) );
  CNIVX1 U3456 ( .A(n256), .Z(n4579) );
  CNIVX1 U3457 ( .A(n4581), .Z(n4580) );
  CNIVX1 U3458 ( .A(n1459), .Z(n4581) );
  CNIVX1 U3459 ( .A(n4583), .Z(n4582) );
  CNIVX1 U3460 ( .A(n1461), .Z(n4583) );
  CNIVX1 U3461 ( .A(n4585), .Z(n4584) );
  CNIVX1 U3462 ( .A(n1463), .Z(n4585) );
  CNIVX1 U3463 ( .A(n4587), .Z(n4586) );
  CNIVX1 U3464 ( .A(n1465), .Z(n4587) );
  CNIVX1 U3465 ( .A(n4589), .Z(n4588) );
  CNIVX1 U3466 ( .A(n1467), .Z(n4589) );
  CNIVX1 U3467 ( .A(n4591), .Z(n4590) );
  CNIVX1 U3468 ( .A(n1469), .Z(n4591) );
  CNIVX1 U3469 ( .A(n4593), .Z(n4592) );
  CNIVX1 U3470 ( .A(n1471), .Z(n4593) );
  CNIVX1 U3471 ( .A(n4595), .Z(n4594) );
  CNIVX1 U3472 ( .A(n1473), .Z(n4595) );
  CNIVX1 U3473 ( .A(n4597), .Z(n4596) );
  CNIVX1 U3474 ( .A(n1475), .Z(n4597) );
  CNIVX1 U3475 ( .A(n4599), .Z(n4598) );
  CNIVX1 U3476 ( .A(n1477), .Z(n4599) );
  CNIVX1 U3477 ( .A(n4601), .Z(n4600) );
  CNIVX1 U3478 ( .A(n1479), .Z(n4601) );
  CNIVX1 U3479 ( .A(n4603), .Z(n4602) );
  CNIVX1 U3480 ( .A(n1457), .Z(n4603) );
  CNIVX1 U3481 ( .A(n4605), .Z(n4604) );
  CNIVX1 U3482 ( .A(n1455), .Z(n4605) );
  CNIVX1 U3483 ( .A(n4607), .Z(n4606) );
  CNIVX1 U3484 ( .A(n1453), .Z(n4607) );
  CNIVX1 U3485 ( .A(n4609), .Z(n4608) );
  CNIVX1 U3486 ( .A(n1451), .Z(n4609) );
  CNIVX1 U3487 ( .A(n4611), .Z(n4610) );
  CNIVX1 U3488 ( .A(n1449), .Z(n4611) );
  CNIVX1 U3489 ( .A(n4613), .Z(n4612) );
  CNIVX1 U3490 ( .A(n1447), .Z(n4613) );
  CNIVX1 U3491 ( .A(n4615), .Z(n4614) );
  CNIVX1 U3492 ( .A(n1445), .Z(n4615) );
  CNIVX1 U3493 ( .A(n4617), .Z(n4616) );
  CNIVX1 U3494 ( .A(n1443), .Z(n4617) );
  CNIVX1 U3495 ( .A(n4619), .Z(n4618) );
  CNIVX1 U3496 ( .A(n1441), .Z(n4619) );
  CNIVX1 U3497 ( .A(n4621), .Z(n4620) );
  CNIVX1 U3498 ( .A(n1439), .Z(n4621) );
  CNIVX1 U3499 ( .A(n4623), .Z(n4622) );
  CNIVX1 U3500 ( .A(n1437), .Z(n4623) );
  CNIVX1 U3501 ( .A(n4625), .Z(n4624) );
  CNIVX1 U3502 ( .A(n1435), .Z(n4625) );
  CNIVX1 U3503 ( .A(n4627), .Z(n4626) );
  CNIVX1 U3504 ( .A(n1433), .Z(n4627) );
  CNIVX1 U3505 ( .A(n4629), .Z(n4628) );
  CNIVX1 U3506 ( .A(n1431), .Z(n4629) );
  CNIVX1 U3507 ( .A(n4631), .Z(n4630) );
  CNIVX1 U3508 ( .A(n1429), .Z(n4631) );
  CNIVX1 U3509 ( .A(n4633), .Z(n4632) );
  CNIVX1 U3510 ( .A(n1460), .Z(n4633) );
  CNIVX1 U3511 ( .A(n4635), .Z(n4634) );
  CNIVX1 U3512 ( .A(n1462), .Z(n4635) );
  CNIVX1 U3513 ( .A(n4637), .Z(n4636) );
  CNIVX1 U3514 ( .A(n1464), .Z(n4637) );
  CNIVX1 U3515 ( .A(n4639), .Z(n4638) );
  CNIVX1 U3516 ( .A(n1466), .Z(n4639) );
  CNIVX1 U3517 ( .A(n4641), .Z(n4640) );
  CNIVX1 U3518 ( .A(n1468), .Z(n4641) );
  CNIVX1 U3519 ( .A(n4643), .Z(n4642) );
  CNIVX1 U3520 ( .A(n1470), .Z(n4643) );
  CNIVX1 U3521 ( .A(n4645), .Z(n4644) );
  CNIVX1 U3522 ( .A(n1472), .Z(n4645) );
  CNIVX1 U3523 ( .A(n4647), .Z(n4646) );
  CNIVX1 U3524 ( .A(n1474), .Z(n4647) );
  CNIVX1 U3525 ( .A(n4649), .Z(n4648) );
  CNIVX1 U3526 ( .A(n1476), .Z(n4649) );
  CNIVX1 U3527 ( .A(n4651), .Z(n4650) );
  CNIVX1 U3528 ( .A(n1478), .Z(n4651) );
  CNIVX1 U3529 ( .A(n4653), .Z(n4652) );
  CNIVX1 U3530 ( .A(n1480), .Z(n4653) );
  CNIVX1 U3531 ( .A(n4655), .Z(n4654) );
  CNIVX1 U3532 ( .A(n1458), .Z(n4655) );
  CNIVX1 U3533 ( .A(n4657), .Z(n4656) );
  CNIVX1 U3534 ( .A(n1456), .Z(n4657) );
  CNIVX1 U3535 ( .A(n4659), .Z(n4658) );
  CNIVX1 U3536 ( .A(n1454), .Z(n4659) );
  CNIVX1 U3537 ( .A(n4661), .Z(n4660) );
  CNIVX1 U3538 ( .A(n1452), .Z(n4661) );
  CNIVX1 U3539 ( .A(n4663), .Z(n4662) );
  CNIVX1 U3540 ( .A(n1450), .Z(n4663) );
  CNIVX1 U3541 ( .A(n4665), .Z(n4664) );
  CNIVX1 U3542 ( .A(n1448), .Z(n4665) );
  CNIVX1 U3543 ( .A(n4667), .Z(n4666) );
  CNIVX1 U3544 ( .A(n1446), .Z(n4667) );
  CNIVX1 U3545 ( .A(n4669), .Z(n4668) );
  CNIVX1 U3546 ( .A(n1444), .Z(n4669) );
  CNIVX1 U3547 ( .A(n4671), .Z(n4670) );
  CNIVX1 U3548 ( .A(n1442), .Z(n4671) );
  CNIVX1 U3549 ( .A(n4673), .Z(n4672) );
  CNIVX1 U3550 ( .A(n1440), .Z(n4673) );
  CNIVX1 U3551 ( .A(n4675), .Z(n4674) );
  CNIVX1 U3552 ( .A(n1438), .Z(n4675) );
  CNIVX1 U3553 ( .A(n4677), .Z(n4676) );
  CNIVX1 U3554 ( .A(n1436), .Z(n4677) );
  CNIVX1 U3555 ( .A(n4679), .Z(n4678) );
  CNIVX1 U3556 ( .A(n1434), .Z(n4679) );
  CNIVX1 U3557 ( .A(n4681), .Z(n4680) );
  CNIVX1 U3558 ( .A(n1432), .Z(n4681) );
  CNIVX1 U3559 ( .A(n4683), .Z(n4682) );
  CNIVX1 U3560 ( .A(n1430), .Z(n4683) );
  CNIVX1 U3561 ( .A(n4685), .Z(n4684) );
  CNIVX1 U3562 ( .A(n1428), .Z(n4685) );
  CNIVX1 U3563 ( .A(n1560), .Z(n4686) );
  CNIVX1 U3564 ( .A(n4134), .Z(n4687) );
  CENXL U3565 ( .A(opera2[60]), .B(n4478), .Z(n4135) );
  COND3XL U3566 ( .A(n3085), .B(n3103), .C(n3495), .D(n3496), .Z(n254) );
  CNIVX1 U3567 ( .A(n4689), .Z(n4688) );
  CNIVX1 U3568 ( .A(n254), .Z(n4689) );
  CNR2IXL U3569 ( .B(opera1_copydiv[31]), .A(n4481), .Z(n3734) );
  CND2XL U3570 ( .A(n3106), .B(n3729), .Z(n3730) );
  CDLY1XL U3571 ( .A(opera1[30]), .Z(n4690) );
  CND4XL U3572 ( .A(n4144), .B(n4145), .C(n4146), .D(n4147), .Z(n1558) );
  CNIVX1 U3573 ( .A(n4692), .Z(n4691) );
  CNIVX1 U3574 ( .A(n1558), .Z(n4692) );
  CNIVX1 U3575 ( .A(n4696), .Z(n4693) );
  CNIVX1 U3576 ( .A(n4695), .Z(n4694) );
  CNIVX1 U3577 ( .A(n4698), .Z(n4695) );
  CNIVX1 U3578 ( .A(n1657), .Z(n4696) );
  CNIVX1 U3579 ( .A(opera1[28]), .Z(n4697) );
  CNIVX1 U3580 ( .A(opera1[29]), .Z(n4698) );
  CNIVX1 U3581 ( .A(n4701), .Z(n4699) );
  CNIVX1 U3582 ( .A(n4703), .Z(n4700) );
  CNIVX1 U3583 ( .A(n1659), .Z(n4701) );
  CNIVX1 U3584 ( .A(opera1[26]), .Z(n4702) );
  CNIVX1 U3585 ( .A(opera1[27]), .Z(n4703) );
  CNIVX1 U3586 ( .A(n1494), .Z(n4704) );
  CNIVX1 U3587 ( .A(n1500), .Z(n4705) );
  CNIVX1 U3588 ( .A(n1498), .Z(n4706) );
  CNIVX1 U3589 ( .A(n1496), .Z(n4707) );
  CNIVX1 U3590 ( .A(n1621), .Z(n4709) );
  COND3X2 U3591 ( .A(n3759), .B(n3276), .C(n3760), .D(n3761), .Z(n1621) );
  CNIVX1 U3592 ( .A(opera2[62]), .Z(n4710) );
  CNR2XL U3593 ( .A(n4136), .B(n4142), .Z(n3765) );
  CEOXL U3594 ( .A(n4710), .B(n4479), .Z(n3767) );
  CNIVXL U3595 ( .A(n250), .Z(n4713) );
  CNIVX1 U3596 ( .A(n4712), .Z(n4711) );
  CNIVX1 U3597 ( .A(n4713), .Z(n4712) );
  COND3X2 U3598 ( .A(n3386), .B(n4477), .C(n3516), .D(n3517), .Z(n250) );
  CNIVX1 U3599 ( .A(n4715), .Z(n4714) );
  CNIVX1 U3600 ( .A(n1629), .Z(n4715) );
  CNIVX1 U3601 ( .A(n4717), .Z(n4716) );
  CNIVXL U3602 ( .A(opera1[21]), .Z(n4817) );
  CNIVX1 U3603 ( .A(n247), .Z(n4717) );
  COND3X2 U3604 ( .A(n3398), .B(n4477), .C(n3530), .D(n3531), .Z(n247) );
  CNIVX1 U3605 ( .A(n4719), .Z(n4718) );
  CNIVX1 U3606 ( .A(n1666), .Z(n4719) );
  CIVXL U3607 ( .A(opera1_copydiv[22]), .Z(n3400) );
  CNIVX1 U3608 ( .A(n4721), .Z(n4720) );
  CNIVX1 U3609 ( .A(n4723), .Z(n4721) );
  CNIVX1 U3610 ( .A(n1664), .Z(n4722) );
  CNIVX1 U3611 ( .A(opera1[22]), .Z(n4723) );
  CNIVX1 U3612 ( .A(n4725), .Z(n4724) );
  CNIVX1 U3613 ( .A(n1662), .Z(n4725) );
  CNIVX1 U3614 ( .A(n246), .Z(n4726) );
  COND3X2 U3615 ( .A(n3402), .B(n4477), .C(n3089), .D(n3536), .Z(n246) );
  CNIVX1 U3616 ( .A(n4729), .Z(n4727) );
  COND3X2 U3617 ( .A(n3403), .B(n4477), .C(n3520), .D(n3521), .Z(n249) );
  CNIVX1 U3618 ( .A(n4731), .Z(n4728) );
  CNIVX1 U3619 ( .A(n4730), .Z(n4729) );
  CNIVX1 U3620 ( .A(n249), .Z(n4730) );
  CNIVX1 U3621 ( .A(opera1[24]), .Z(n4731) );
  COND3X2 U3622 ( .A(n3404), .B(n4477), .C(n3526), .D(n3527), .Z(n248) );
  CNIVX1 U3623 ( .A(n4733), .Z(n4732) );
  CNIVX1 U3624 ( .A(n248), .Z(n4733) );
  CNIVX1 U3625 ( .A(n4736), .Z(n4734) );
  CNIVX1 U3626 ( .A(n4738), .Z(n4735) );
  CNIVX1 U3627 ( .A(n4737), .Z(n4736) );
  CNIVX1 U3628 ( .A(n4814), .Z(n4737) );
  CNIVX1 U3629 ( .A(n245), .Z(n4738) );
  CNIVXL U3630 ( .A(n244), .Z(n4740) );
  COND3X2 U3631 ( .A(n3406), .B(n4477), .C(n3547), .D(n3548), .Z(n244) );
  CNIVX1 U3632 ( .A(n4740), .Z(n4739) );
  CNIVX1 U3633 ( .A(n4742), .Z(n4741) );
  CNIVX1 U3634 ( .A(n1626), .Z(n4742) );
  CNIVX1 U3635 ( .A(n4744), .Z(n4743) );
  CNIVX1 U3636 ( .A(n1634), .Z(n4744) );
  CNIVX1 U3637 ( .A(n4746), .Z(n4745) );
  CNIVX1 U3638 ( .A(n1642), .Z(n4746) );
  CNIVX1 U3639 ( .A(n4748), .Z(n4747) );
  CNIVX1 U3640 ( .A(n1648), .Z(n4748) );
  CNIVX1 U3641 ( .A(n4750), .Z(n4749) );
  CNIVX1 U3642 ( .A(n1650), .Z(n4750) );
  CNIVX1 U3643 ( .A(n4752), .Z(n4751) );
  CNIVX1 U3644 ( .A(n1640), .Z(n4752) );
  CNIVX1 U3645 ( .A(n4754), .Z(n4753) );
  CNIVX1 U3646 ( .A(n1638), .Z(n4754) );
  CNIVX1 U3647 ( .A(n4756), .Z(n4755) );
  CNIVX1 U3648 ( .A(n1636), .Z(n4756) );
  CNIVX1 U3649 ( .A(n4758), .Z(n4757) );
  CNIVX1 U3650 ( .A(n1628), .Z(n4758) );
  CNIVX1 U3651 ( .A(n4760), .Z(n4759) );
  CNIVX1 U3652 ( .A(n1632), .Z(n4760) );
  CNIVX1 U3653 ( .A(n4762), .Z(n4761) );
  CNIVX1 U3654 ( .A(n1630), .Z(n4762) );
  CNIVX1 U3655 ( .A(n4764), .Z(n4763) );
  CNIVX1 U3656 ( .A(n1646), .Z(n4764) );
  CNIVX1 U3657 ( .A(n4766), .Z(n4765) );
  CNIVX1 U3658 ( .A(n1644), .Z(n4766) );
  CNIVX1 U3659 ( .A(n4768), .Z(n4767) );
  CNIVX1 U3660 ( .A(n1627), .Z(n4768) );
  CNIVX1 U3661 ( .A(n4770), .Z(n4769) );
  CNIVX1 U3662 ( .A(n1649), .Z(n4770) );
  CNIVX1 U3663 ( .A(n4772), .Z(n4771) );
  CNIVX1 U3664 ( .A(n1639), .Z(n4772) );
  CNIVX1 U3665 ( .A(n4774), .Z(n4773) );
  CNIVX1 U3666 ( .A(n1647), .Z(n4774) );
  CNIVX1 U3667 ( .A(n4776), .Z(n4775) );
  CNIVX1 U3668 ( .A(n1631), .Z(n4776) );
  CNIVX1 U3669 ( .A(n4778), .Z(n4777) );
  CNIVX1 U3670 ( .A(n1643), .Z(n4778) );
  CNIVX1 U3671 ( .A(n4780), .Z(n4779) );
  CNIVX1 U3672 ( .A(n1633), .Z(n4780) );
  CNIVX1 U3673 ( .A(n4782), .Z(n4781) );
  CNIVX1 U3674 ( .A(n1645), .Z(n4782) );
  CNIVX1 U3675 ( .A(n4784), .Z(n4783) );
  CNIVX1 U3676 ( .A(n1641), .Z(n4784) );
  CNIVX1 U3677 ( .A(n4786), .Z(n4785) );
  CNIVX1 U3678 ( .A(n1635), .Z(n4786) );
  CNIVX1 U3679 ( .A(n4788), .Z(n4787) );
  CNIVX1 U3680 ( .A(n1637), .Z(n4788) );
  CIVXL U3681 ( .A(i[1]), .Z(n3440) );
  CNIVX1 U3682 ( .A(n1624), .Z(n4789) );
  CNIVX1 U3683 ( .A(n4791), .Z(n4790) );
  CNIVX1 U3684 ( .A(n1653), .Z(n4791) );
  CNIVX2 U3685 ( .A(n1625), .Z(n4792) );
  CNIVX1 U3686 ( .A(n4794), .Z(n4793) );
  CNIVX1 U3687 ( .A(n1564), .Z(n4795) );
  CNIVX1 U3688 ( .A(n4108), .Z(n4796) );
  CENXL U3689 ( .A(opera2[56]), .B(n4478), .Z(n4109) );
  CNIVX1 U3690 ( .A(n1568), .Z(n4797) );
  CNIVX1 U3691 ( .A(n4082), .Z(n4798) );
  CENXL U3692 ( .A(opera2[52]), .B(n4478), .Z(n4083) );
  COND3X2 U3693 ( .A(n3746), .B(n3439), .C(n3750), .D(n3749), .Z(n1623) );
  CNIVX1 U3694 ( .A(n4800), .Z(n4799) );
  CNIVX1 U3695 ( .A(n1652), .Z(n4800) );
  CNIVX1 U3696 ( .A(n4804), .Z(n4801) );
  CNIVX1 U3697 ( .A(n4120), .Z(n4802) );
  CNIVX1 U3698 ( .A(n4121), .Z(n4803) );
  CNIVX1 U3699 ( .A(n1562), .Z(n4804) );
  CEOXL U3700 ( .A(opera2[58]), .B(n4478), .Z(n4122) );
  CNIVX1 U3701 ( .A(n4808), .Z(n4805) );
  CNIVX1 U3702 ( .A(n4094), .Z(n4806) );
  CNIVX1 U3703 ( .A(n4095), .Z(n4807) );
  CNIVX1 U3704 ( .A(n1566), .Z(n4808) );
  CEOXL U3705 ( .A(opera2[54]), .B(n4478), .Z(n4096) );
  COND11XL U3706 ( .A(n3741), .B(n3360), .C(n3283), .D(n3742), .Z(n1651) );
  CNIVX1 U3707 ( .A(n1651), .Z(n4809) );
  CNIVX1 U3708 ( .A(n4811), .Z(n4810) );
  CNIVX1 U3709 ( .A(n1661), .Z(n4811) );
  CNIVX1 U3710 ( .A(n4816), .Z(n4813) );
  CNIVX1 U3711 ( .A(opera1[20]), .Z(n4814) );
  CNIVX1 U3712 ( .A(n3146), .Z(n4815) );
  CNIVX1 U3713 ( .A(n1665), .Z(n4816) );
  CNIVX1 U3714 ( .A(n4821), .Z(n4818) );
  CNIVX1 U3715 ( .A(n4820), .Z(n4819) );
  CNIVX1 U3716 ( .A(n1663), .Z(n4820) );
  CNIVX1 U3717 ( .A(opera1[23]), .Z(n4821) );
  CNIVX1 U3718 ( .A(n1508), .Z(n4822) );
  CNIVX1 U3719 ( .A(n1506), .Z(n4823) );
  CNIVX1 U3720 ( .A(n1504), .Z(n4824) );
  CNIVX1 U3721 ( .A(n1502), .Z(n4825) );
  CNIVX1 U3722 ( .A(n1510), .Z(n4826) );
  CIVDX1 U3723 ( .A(nest[1]), .Z1(n4829) );
  CNIVX1 U3724 ( .A(n4829), .Z(n4828) );
  CNIVX1 U3725 ( .A(n4831), .Z(n4830) );
  CNIVX1 U3726 ( .A(n4832), .Z(n4831) );
  CNIVX1 U3727 ( .A(n243), .Z(n4832) );
  CNIVX1 U3728 ( .A(n4834), .Z(n4833) );
  CNIVX1 U3729 ( .A(n4835), .Z(n4834) );
  CNIVX1 U3730 ( .A(n239), .Z(n4835) );
  CIVXL U3731 ( .A(opera1_copydiv[14]), .Z(n3443) );
  CNIVX1 U3732 ( .A(n4837), .Z(n4836) );
  CNIVX1 U3733 ( .A(n4878), .Z(n4837) );
  CNIVX1 U3734 ( .A(n1672), .Z(n4838) );
  CNIVX1 U3735 ( .A(n4840), .Z(n4839) );
  CNIVX1 U3736 ( .A(n1670), .Z(n4840) );
  COND4CXL U3737 ( .A(n3117), .B(n3134), .C(n3692), .D(n3693), .Z(n3691) );
  CIVXL U3738 ( .A(opera1_copydiv[18]), .Z(n3445) );
  CNIVX1 U3739 ( .A(n4842), .Z(n4841) );
  CNIVX1 U3740 ( .A(n4872), .Z(n4842) );
  CNIVX1 U3741 ( .A(n1668), .Z(n4843) );
  COND3XL U3742 ( .A(n3446), .B(n4477), .C(n3088), .D(n3557), .Z(n242) );
  CNIVX1 U3743 ( .A(n4845), .Z(n4844) );
  CNIVX1 U3744 ( .A(n242), .Z(n4845) );
  COND3XL U3745 ( .A(n3447), .B(n4477), .C(n3087), .D(n3577), .Z(n238) );
  CNIVX1 U3746 ( .A(n4847), .Z(n4846) );
  CNIVX1 U3747 ( .A(n238), .Z(n4847) );
  CNIVX2 U3748 ( .A(n241), .Z(n4848) );
  CDLY1XL U3749 ( .A(opera1[16]), .Z(n4865) );
  COND3X2 U3750 ( .A(n3449), .B(n4477), .C(n3567), .D(n3568), .Z(n240) );
  CNIVX1 U3751 ( .A(n240), .Z(n4849) );
  CNIVX1 U3752 ( .A(n1572), .Z(n4850) );
  CNIVX1 U3753 ( .A(n4056), .Z(n4851) );
  CENXL U3754 ( .A(opera2[48]), .B(n4478), .Z(n4057) );
  CNIVX1 U3755 ( .A(n4855), .Z(n4852) );
  CNIVX1 U3756 ( .A(n4068), .Z(n4853) );
  CNIVX1 U3757 ( .A(n4069), .Z(n4854) );
  CNIVX1 U3758 ( .A(n1570), .Z(n4855) );
  CEOXL U3759 ( .A(opera2[50]), .B(n4478), .Z(n4070) );
  CNIVX1 U3760 ( .A(n4859), .Z(n4856) );
  CNIVX1 U3761 ( .A(n4042), .Z(n4857) );
  CNIVX1 U3762 ( .A(n4043), .Z(n4858) );
  CNIVX1 U3763 ( .A(n1574), .Z(n4859) );
  CEOXL U3764 ( .A(opera2[46]), .B(n4478), .Z(n4044) );
  CNIVX1 U3765 ( .A(n4861), .Z(n4860) );
  CNIVX1 U3766 ( .A(n1673), .Z(n4861) );
  CNIVX1 U3767 ( .A(n3154), .Z(n4862) );
  CNIVX1 U3768 ( .A(opera1[13]), .Z(n4863) );
  CNIVX1 U3769 ( .A(n4867), .Z(n4864) );
  CNIVX1 U3770 ( .A(n3150), .Z(n4866) );
  CNIVX1 U3771 ( .A(n1669), .Z(n4867) );
  CNIVX1 U3772 ( .A(opera1[17]), .Z(n4868) );
  CNIVX1 U3773 ( .A(n4871), .Z(n4869) );
  CNIVX1 U3774 ( .A(n4873), .Z(n4870) );
  CNIVX1 U3775 ( .A(n1667), .Z(n4871) );
  CNIVX1 U3776 ( .A(opera1[18]), .Z(n4872) );
  CNIVX1 U3777 ( .A(opera1[19]), .Z(n4873) );
  CNIVX1 U3778 ( .A(n4877), .Z(n4874) );
  CNIVX1 U3779 ( .A(n4876), .Z(n4875) );
  CNIVX1 U3780 ( .A(n4879), .Z(n4876) );
  CNIVX1 U3781 ( .A(n1671), .Z(n4877) );
  CNIVX1 U3782 ( .A(opera1[14]), .Z(n4878) );
  CNIVX1 U3783 ( .A(opera1[15]), .Z(n4879) );
  CNIVX1 U3784 ( .A(n1518), .Z(n4880) );
  CNIVX1 U3785 ( .A(n1516), .Z(n4881) );
  CNIVX1 U3786 ( .A(n1514), .Z(n4882) );
  CNIVX1 U3787 ( .A(n1512), .Z(n4883) );
  CNIVX1 U3788 ( .A(n4885), .Z(n4884) );
  CNIVX1 U3789 ( .A(n4886), .Z(n4885) );
  CNIVX1 U3790 ( .A(n237), .Z(n4886) );
  CNIVX1 U3791 ( .A(n4888), .Z(n4887) );
  CNIVX1 U3792 ( .A(n4889), .Z(n4888) );
  CNIVX1 U3793 ( .A(n235), .Z(n4889) );
  CNIVX1 U3794 ( .A(n4891), .Z(n4890) );
  CNIVX1 U3795 ( .A(n4892), .Z(n4891) );
  CNIVX1 U3796 ( .A(n231), .Z(n4892) );
  CNIVX1 U3797 ( .A(n4894), .Z(n4893) );
  CNIVX1 U3798 ( .A(n1678), .Z(n4894) );
  CIVXL U3799 ( .A(opera1_copydiv[10]), .Z(n3458) );
  CNIVX1 U3800 ( .A(n4896), .Z(n4895) );
  CNIVX1 U3801 ( .A(n4930), .Z(n4896) );
  CNIVX1 U3802 ( .A(n1676), .Z(n4897) );
  CNIVX1 U3803 ( .A(n4901), .Z(n4898) );
  CNIVX1 U3804 ( .A(n4900), .Z(n4899) );
  CNIVX1 U3805 ( .A(n4902), .Z(n4900) );
  CNIVX1 U3806 ( .A(n1674), .Z(n4901) );
  CNIVX1 U3807 ( .A(opera1[12]), .Z(n4902) );
  COND3XL U3808 ( .A(n3460), .B(n4477), .C(n3086), .D(n3597), .Z(n234) );
  CNIVX1 U3809 ( .A(n4904), .Z(n4903) );
  CNIVX1 U3810 ( .A(n234), .Z(n4904) );
  CNIVXL U3811 ( .A(n236), .Z(n4906) );
  COND3X2 U3812 ( .A(n3461), .B(n4477), .C(n3587), .D(n3588), .Z(n236) );
  CNIVX1 U3813 ( .A(n4906), .Z(n4905) );
  CNIVX2 U3814 ( .A(n233), .Z(n4907) );
  CDLY1XL U3815 ( .A(opera1[8]), .Z(n4920) );
  COND3X2 U3816 ( .A(n3463), .B(n4477), .C(n3607), .D(n3608), .Z(n232) );
  CNIVX1 U3817 ( .A(n232), .Z(n4908) );
  CNIVX1 U3818 ( .A(n1576), .Z(n4909) );
  CNIVX1 U3819 ( .A(n4030), .Z(n4910) );
  CENXL U3820 ( .A(opera2[44]), .B(n4478), .Z(n4031) );
  CNIVX1 U3821 ( .A(n1580), .Z(n4911) );
  CNIVX1 U3822 ( .A(n4004), .Z(n4912) );
  CENXL U3823 ( .A(opera2[40]), .B(n4478), .Z(n4005) );
  CNIVX1 U3824 ( .A(n4916), .Z(n4913) );
  CNIVX1 U3825 ( .A(n4016), .Z(n4914) );
  CNIVX1 U3826 ( .A(n4017), .Z(n4915) );
  CNIVX1 U3827 ( .A(n1578), .Z(n4916) );
  CEOXL U3828 ( .A(opera2[42]), .B(n4478), .Z(n4018) );
  CNIVX1 U3829 ( .A(n4918), .Z(n4917) );
  CNIVX1 U3830 ( .A(n1677), .Z(n4918) );
  CNIVX1 U3831 ( .A(n3158), .Z(n4919) );
  CNIVX1 U3832 ( .A(opera1[9]), .Z(n4921) );
  CNIVX1 U3833 ( .A(n4925), .Z(n4922) );
  CNIVX1 U3834 ( .A(n4924), .Z(n4923) );
  CNIVX1 U3835 ( .A(n4926), .Z(n4924) );
  CNIVX1 U3836 ( .A(n1679), .Z(n4925) );
  CNIVX1 U3837 ( .A(opera1[7]), .Z(n4926) );
  CNIVX1 U3838 ( .A(n4929), .Z(n4927) );
  CNIVX1 U3839 ( .A(n4931), .Z(n4928) );
  CNIVX1 U3840 ( .A(n1675), .Z(n4929) );
  CNIVX1 U3841 ( .A(opera1[10]), .Z(n4930) );
  CNIVX1 U3842 ( .A(opera1[11]), .Z(n4931) );
  CNIVX1 U3843 ( .A(n1520), .Z(n4932) );
  CNIVX1 U3844 ( .A(n1524), .Z(n4933) );
  COND3X2 U3845 ( .A(n3948), .B(n4143), .C(n4210), .D(n4211), .Z(n1522) );
  CNIVX1 U3846 ( .A(n1526), .Z(n4934) );
  CIVXL U3847 ( .A(opera1_copydiv[6]), .Z(n3456) );
  CNIVX1 U3848 ( .A(n4936), .Z(n4935) );
  CNIVX1 U3849 ( .A(n4938), .Z(n4936) );
  CNIVX1 U3850 ( .A(n1680), .Z(n4937) );
  CNIVX1 U3851 ( .A(opera1[6]), .Z(n4938) );
  CNIVX1 U3852 ( .A(n4940), .Z(n4939) );
  CNIVX1 U3853 ( .A(n4941), .Z(n4940) );
  CNIVX1 U3854 ( .A(n227), .Z(n4941) );
  CNIVX1 U3855 ( .A(n4945), .Z(n4942) );
  CNIVX1 U3856 ( .A(n4944), .Z(n4943) );
  CNIVX1 U3857 ( .A(n4946), .Z(n4944) );
  CNIVX1 U3858 ( .A(n1684), .Z(n4945) );
  CNIVX1 U3859 ( .A(opera1[2]), .Z(n4946) );
  COND4CXL U3860 ( .A(n3129), .B(n3657), .C(n3659), .D(n3660), .Z(n3658) );
  CNIVX1 U3861 ( .A(n4948), .Z(n4947) );
  CNIVX1 U3862 ( .A(n1682), .Z(n4948) );
  CNIVXL U3863 ( .A(n230), .Z(n4949) );
  COND3X2 U3864 ( .A(n3470), .B(n4477), .C(n3100), .D(n3617), .Z(n230) );
  CNIVX1 U3865 ( .A(n3621), .Z(n4950) );
  CNIVX1 U3866 ( .A(n4953), .Z(n4951) );
  CNIVX1 U3867 ( .A(n4968), .Z(n4952) );
  CNIVX1 U3868 ( .A(n229), .Z(n4953) );
  CDLY1XL U3869 ( .A(n228), .Z(n4954) );
  COND3XL U3870 ( .A(n3472), .B(n4477), .C(n3627), .D(n3628), .Z(n228) );
  COND3X2 U3871 ( .A(n3473), .B(n4477), .C(n3637), .D(n3638), .Z(n226) );
  CNIVX1 U3872 ( .A(n226), .Z(n4955) );
  CIVX3 U3873 ( .A(opera1_copydiv[0]), .Z(n3474) );
  CNIVX1 U3874 ( .A(n1686), .Z(n4956) );
  CNIVXL U3875 ( .A(opera1[31]), .Z(n4986) );
  CNIVX1 U3876 ( .A(n4960), .Z(n4957) );
  CNIVX1 U3877 ( .A(n3962), .Z(n4958) );
  CNIVX1 U3878 ( .A(n3963), .Z(n4959) );
  CNIVX1 U3879 ( .A(n1586), .Z(n4960) );
  CEOXL U3880 ( .A(opera2[34]), .B(n4478), .Z(n3964) );
  CNIVX1 U3881 ( .A(n4964), .Z(n4961) );
  CNIVX1 U3882 ( .A(n3990), .Z(n4962) );
  CNIVX1 U3883 ( .A(n3991), .Z(n4963) );
  CNIVX1 U3884 ( .A(n1582), .Z(n4964) );
  CEOXL U3885 ( .A(opera2[38]), .B(n4478), .Z(n3992) );
  CNIVX1 U3886 ( .A(n4966), .Z(n4965) );
  CNIVX1 U3887 ( .A(n1681), .Z(n4966) );
  CNIVX1 U3888 ( .A(n3161), .Z(n4967) );
  CNIVX1 U3889 ( .A(opera1[4]), .Z(n4968) );
  CNIVX1 U3890 ( .A(opera1[5]), .Z(n4969) );
  CNIVX1 U3891 ( .A(n4973), .Z(n4970) );
  CNIVX1 U3892 ( .A(n4972), .Z(n4971) );
  CNIVX1 U3893 ( .A(n4974), .Z(n4972) );
  CNIVX1 U3894 ( .A(n1685), .Z(n4973) );
  CNIVX1 U3895 ( .A(opera1[1]), .Z(n4974) );
  CNIVX1 U3896 ( .A(n4976), .Z(n4975) );
  CNIVX1 U3897 ( .A(n1683), .Z(n4976) );
  CNIVX1 U3898 ( .A(opera1[3]), .Z(n4977) );
  CNIVX1 U3899 ( .A(n1528), .Z(n4978) );
  CNIVX1 U3900 ( .A(n1530), .Z(n4979) );
  CNIVX1 U3901 ( .A(n1532), .Z(n4980) );
  CNIVX1 U3902 ( .A(n1534), .Z(n4981) );
  CNIVX1 U3903 ( .A(n1536), .Z(n4982) );
  COND3X2 U3904 ( .A(n4486), .B(n3641), .C(n3642), .D(n3643), .Z(n225) );
  CNIVX1 U3905 ( .A(n4988), .Z(n4983) );
  CNIVX1 U3906 ( .A(n4985), .Z(n4984) );
  CNIVX1 U3907 ( .A(n4987), .Z(n4985) );
  CNIVX1 U3908 ( .A(opera1[0]), .Z(n4987) );
  CNIVX1 U3909 ( .A(n225), .Z(n4988) );
  CANR2XL U3910 ( .A(n4984), .B(n3640), .C(opera1_copy[0]), .D(n4476), .Z(
        n3643) );
  CNIVX1 U3911 ( .A(n4992), .Z(n4989) );
  CNIVX1 U3912 ( .A(n3940), .Z(n4990) );
  CNIVX1 U3913 ( .A(n3941), .Z(n4991) );
  CNIVX1 U3914 ( .A(n1588), .Z(n4992) );
  CEOXL U3915 ( .A(opera2[32]), .B(n4478), .Z(n3946) );
  CNIVX1 U3916 ( .A(n1584), .Z(n4993) );
  CNIVX1 U3917 ( .A(n3978), .Z(n4994) );
  CENXL U3918 ( .A(opera2[36]), .B(n4478), .Z(n3979) );
  CNIVX1 U3919 ( .A(n1538), .Z(n4995) );
  CNIVX1 U3920 ( .A(n1540), .Z(n4996) );
  CNIVX1 U3921 ( .A(n1542), .Z(n4997) );
  CNIVX1 U3922 ( .A(n1544), .Z(n4998) );
  CNIVX1 U3923 ( .A(n224), .Z(n4999) );
  CNR2XL U3924 ( .A(n4476), .B(n4986), .Z(n3545) );
  CNIVX1 U3925 ( .A(n1546), .Z(n5000) );
  CNIVX1 U3926 ( .A(n1550), .Z(n5001) );
  COND3X2 U3927 ( .A(n3763), .B(n4143), .C(n4175), .D(n4176), .Z(n1554) );
  CNIVX1 U3928 ( .A(n1548), .Z(n5002) );
  CNIVX1 U3929 ( .A(n1552), .Z(n5003) );
  CND2IX2 U3930 ( .B(n5008), .A(n5005), .Z(n257) );
  CNIVX1 U3931 ( .A(n257), .Z(n5004) );
  CNIVX1 U3932 ( .A(n5006), .Z(n5005) );
  CNIVX1 U3933 ( .A(nest[2]), .Z(n5006) );
  CDLY1XL U3934 ( .A(nest[0]), .Z(n5007) );
  CDLY2XL U3935 ( .A(start), .Z(n5008) );
  CNIVX1 U3936 ( .A(n5010), .Z(n5009) );
  CNIVX1 U3937 ( .A(result_copy[31]), .Z(n5010) );
  CNIVX1 U3938 ( .A(n1523), .Z(n5011) );
  CNIVX1 U3939 ( .A(n1525), .Z(n5012) );
  CNIVX1 U3940 ( .A(n1527), .Z(n5013) );
  CNIVX1 U3941 ( .A(n1529), .Z(n5014) );
  CNIVX1 U3942 ( .A(n1531), .Z(n5015) );
  CNIVX1 U3943 ( .A(n1533), .Z(n5016) );
  CNIVX1 U3944 ( .A(n1535), .Z(n5017) );
  CNIVX1 U3945 ( .A(n1537), .Z(n5018) );
  CNIVX1 U3946 ( .A(n1539), .Z(n5019) );
  CNIVX1 U3947 ( .A(n1541), .Z(n5020) );
  CNIVX1 U3948 ( .A(n1543), .Z(n5021) );
  CNIVX1 U3949 ( .A(n1545), .Z(n5022) );
  CNIVX1 U3950 ( .A(n5024), .Z(n5023) );
  CNIVX1 U3951 ( .A(n1547), .Z(n5024) );
  CNIVX1 U3952 ( .A(n1549), .Z(n5025) );
  CNIVX1 U3953 ( .A(n5027), .Z(n5026) );
  CNIVX1 U3954 ( .A(n1551), .Z(n5027) );
  CNIVX1 U3955 ( .A(n5029), .Z(n5028) );
  CNIVX1 U3956 ( .A(n1553), .Z(n5029) );
  CNIVX1 U3957 ( .A(n1517), .Z(n5030) );
  CNIVX1 U3958 ( .A(n1519), .Z(n5031) );
  CNIVX1 U3959 ( .A(n1521), .Z(n5032) );
  CNIVX1 U3960 ( .A(n1515), .Z(n5033) );
  CNIVX1 U3961 ( .A(n1611), .Z(n5034) );
  CNIVX1 U3962 ( .A(opera2[8]), .Z(n5035) );
  CDLY1XL U3963 ( .A(opera2[9]), .Z(n5036) );
  CANR2XL U3964 ( .A(n5182), .B(n3822), .C(n5180), .D(n5036), .Z(n3820) );
  CNIVX1 U3965 ( .A(n5038), .Z(n5037) );
  CNIVX1 U3966 ( .A(n5039), .Z(n5038) );
  CNIVX1 U3967 ( .A(n5041), .Z(n5039) );
  CNIVX1 U3968 ( .A(opera2[5]), .Z(n5040) );
  CNIVX1 U3969 ( .A(n1615), .Z(n5041) );
  CANR2XL U3970 ( .A(n5182), .B(n3803), .C(n5180), .D(n5040), .Z(n3801) );
  CNIVX1 U3971 ( .A(n5043), .Z(n5042) );
  CNIVX1 U3972 ( .A(n5044), .Z(n5043) );
  CNIVX1 U3973 ( .A(n5045), .Z(n5044) );
  CNIVX1 U3974 ( .A(n5047), .Z(n5045) );
  CNIVX1 U3975 ( .A(opera2[1]), .Z(n5046) );
  CNIVX1 U3976 ( .A(n1619), .Z(n5047) );
  CANR2XL U3977 ( .A(n3784), .B(n5181), .C(n5180), .D(n5046), .Z(n3781) );
  CNIVX1 U3978 ( .A(n1513), .Z(n5048) );
  CNIVX1 U3979 ( .A(n5050), .Z(n5049) );
  CNIVX1 U3980 ( .A(n5051), .Z(n5050) );
  CNIVX1 U3981 ( .A(n5053), .Z(n5051) );
  CNIVX1 U3982 ( .A(opera2[13]), .Z(n5052) );
  CNIVX1 U3983 ( .A(n1607), .Z(n5053) );
  CANR2XL U3984 ( .A(n3841), .B(n5182), .C(n5180), .D(n5052), .Z(n3839) );
  CNIVX1 U3985 ( .A(n1511), .Z(n5054) );
  CNIVX1 U3986 ( .A(n5056), .Z(n5055) );
  CNIVX1 U3987 ( .A(n5057), .Z(n5056) );
  CNIVX1 U3988 ( .A(n5059), .Z(n5057) );
  CNIVX1 U3989 ( .A(opera2[15]), .Z(n5058) );
  CNIVX1 U3990 ( .A(n1605), .Z(n5059) );
  CANR2XL U3991 ( .A(n5182), .B(n3852), .C(n5180), .D(n5058), .Z(n3850) );
  CNIVX1 U3992 ( .A(n5061), .Z(n5060) );
  CNIVX1 U3993 ( .A(n5062), .Z(n5061) );
  CNIVX1 U3994 ( .A(n5064), .Z(n5062) );
  CNIVX1 U3995 ( .A(opera2[17]), .Z(n5063) );
  CNIVX1 U3996 ( .A(n1603), .Z(n5064) );
  CANR2XL U3997 ( .A(n3862), .B(n5182), .C(n5180), .D(n5063), .Z(n3860) );
  CNIVX1 U3998 ( .A(n5066), .Z(n5065) );
  CNIVX1 U3999 ( .A(n5067), .Z(n5066) );
  CNIVX1 U4000 ( .A(n5069), .Z(n5067) );
  CNIVX1 U4001 ( .A(opera2[19]), .Z(n5068) );
  CNIVX1 U4002 ( .A(n1601), .Z(n5069) );
  CANR2XL U4003 ( .A(n5181), .B(n3873), .C(n5180), .D(n5068), .Z(n3871) );
  CNIVX1 U4004 ( .A(n1509), .Z(n5070) );
  CNIVX1 U4005 ( .A(n5072), .Z(n5071) );
  CNIVX1 U4006 ( .A(n5073), .Z(n5072) );
  CNIVX1 U4007 ( .A(n5075), .Z(n5073) );
  CNIVX1 U4008 ( .A(opera2[21]), .Z(n5074) );
  CNIVX1 U4009 ( .A(n1599), .Z(n5075) );
  CANR2XL U4010 ( .A(n3883), .B(n3778), .C(n5180), .D(n5074), .Z(n3881) );
  CNIVX1 U4011 ( .A(n5077), .Z(n5076) );
  CNIVX1 U4012 ( .A(n5078), .Z(n5077) );
  CNIVX1 U4013 ( .A(n5080), .Z(n5078) );
  CNIVX1 U4014 ( .A(opera2[23]), .Z(n5079) );
  CNIVX1 U4015 ( .A(n1597), .Z(n5080) );
  CANR2XL U4016 ( .A(n5181), .B(n3894), .C(n5180), .D(n5079), .Z(n3892) );
  CNIVX1 U4017 ( .A(n1507), .Z(n5081) );
  CNIVX1 U4018 ( .A(n5083), .Z(n5082) );
  CNIVX1 U4019 ( .A(n5084), .Z(n5083) );
  CNIVX1 U4020 ( .A(n5086), .Z(n5084) );
  CNIVX1 U4021 ( .A(opera2[25]), .Z(n5085) );
  CNIVX1 U4022 ( .A(n1595), .Z(n5086) );
  CANR2XL U4023 ( .A(n3904), .B(n3778), .C(n5180), .D(n5085), .Z(n3902) );
  CNIVX1 U4024 ( .A(n5088), .Z(n5087) );
  CNIVX1 U4025 ( .A(n5089), .Z(n5088) );
  CNIVX1 U4026 ( .A(n5091), .Z(n5089) );
  CNIVX1 U4027 ( .A(opera2[27]), .Z(n5090) );
  CNIVX1 U4028 ( .A(n1593), .Z(n5091) );
  CANR2XL U4029 ( .A(n5181), .B(n3915), .C(n5180), .D(n5090), .Z(n3913) );
  CNIVX1 U4030 ( .A(n1505), .Z(n5092) );
  CNIVX1 U4031 ( .A(n5094), .Z(n5093) );
  CNIVX1 U4032 ( .A(n5095), .Z(n5094) );
  CNIVX1 U4033 ( .A(n5097), .Z(n5095) );
  CNIVX1 U4034 ( .A(opera2[29]), .Z(n5096) );
  CNIVX1 U4035 ( .A(n1591), .Z(n5097) );
  CANR2XL U4036 ( .A(n5181), .B(n3925), .C(n5180), .D(n5096), .Z(n3923) );
  CNIVX1 U4037 ( .A(n1503), .Z(n5098) );
  CNIVX1 U4038 ( .A(n5100), .Z(n5099) );
  CNIVX1 U4039 ( .A(n5102), .Z(n5100) );
  CNIVX1 U4040 ( .A(opera2[31]), .Z(n5101) );
  CNIVX1 U4041 ( .A(n1589), .Z(n5102) );
  CNIVX1 U4042 ( .A(n1501), .Z(n5103) );
  CNIVX1 U4043 ( .A(n1499), .Z(n5104) );
  CNIVX1 U4044 ( .A(n1497), .Z(n5105) );
  CNIVX1 U4045 ( .A(n1495), .Z(n5106) );
  CNIVX1 U4046 ( .A(n1493), .Z(n5107) );
  CNIVX1 U4047 ( .A(n1557), .Z(n5108) );
  CNIVX1 U4048 ( .A(n5111), .Z(n5109) );
  CNIVX1 U4049 ( .A(n3953), .Z(n5110) );
  CENXL U4050 ( .A(opera2[33]), .B(n4479), .Z(n3956) );
  CNIVX1 U4051 ( .A(n1587), .Z(n5111) );
  CNIVX1 U4052 ( .A(opera2[35]), .Z(n5112) );
  CNIVX1 U4053 ( .A(n3971), .Z(n5113) );
  CNIVX1 U4054 ( .A(n1585), .Z(n5114) );
  CENXL U4055 ( .A(n5112), .B(n4478), .Z(n3972) );
  CNIVX1 U4056 ( .A(n5117), .Z(n5115) );
  CNIVX1 U4057 ( .A(n3985), .Z(n5116) );
  CENXL U4058 ( .A(opera2[37]), .B(n4479), .Z(n3986) );
  CNIVX1 U4059 ( .A(n1583), .Z(n5117) );
  CNIVX1 U4060 ( .A(n5119), .Z(n5118) );
  CNIVX1 U4061 ( .A(n5120), .Z(n5119) );
  CENXL U4062 ( .A(opera2[39]), .B(n4478), .Z(n3999) );
  CNIVX1 U4063 ( .A(n1581), .Z(n5120) );
  CNIVX1 U4064 ( .A(n5123), .Z(n5121) );
  CNIVX1 U4065 ( .A(n4011), .Z(n5122) );
  CENXL U4066 ( .A(opera2[41]), .B(n4479), .Z(n4012) );
  CNIVX1 U4067 ( .A(n1579), .Z(n5123) );
  CNIVX1 U4068 ( .A(n5126), .Z(n5124) );
  CNIVX1 U4069 ( .A(n4024), .Z(n5125) );
  CNIVX1 U4070 ( .A(n5127), .Z(n5126) );
  CNIVX1 U4071 ( .A(n1577), .Z(n5127) );
  CNIVX1 U4072 ( .A(n5130), .Z(n5128) );
  CNIVX1 U4073 ( .A(n4037), .Z(n5129) );
  CENXL U4074 ( .A(opera2[45]), .B(n4479), .Z(n4038) );
  CNIVX1 U4075 ( .A(n1575), .Z(n5130) );
  CNIVX1 U4076 ( .A(n5132), .Z(n5131) );
  CNIVX1 U4077 ( .A(n5133), .Z(n5132) );
  CENXL U4078 ( .A(opera2[47]), .B(n4478), .Z(n4051) );
  CNIVX1 U4079 ( .A(n1573), .Z(n5133) );
  CNIVX1 U4080 ( .A(n5136), .Z(n5134) );
  CNIVX1 U4081 ( .A(n4063), .Z(n5135) );
  CENXL U4082 ( .A(opera2[49]), .B(n4479), .Z(n4064) );
  CNIVX1 U4083 ( .A(n1571), .Z(n5136) );
  CNIVX1 U4084 ( .A(n5138), .Z(n5137) );
  CNIVX1 U4085 ( .A(n5139), .Z(n5138) );
  CENXL U4086 ( .A(opera2[51]), .B(n4478), .Z(n4077) );
  CNIVX1 U4087 ( .A(n1569), .Z(n5139) );
  CNIVX1 U4088 ( .A(n5142), .Z(n5140) );
  CNIVX1 U4089 ( .A(opera2[53]), .Z(n5141) );
  CNIVX1 U4090 ( .A(n1567), .Z(n5142) );
  CNIVX1 U4091 ( .A(n5145), .Z(n5143) );
  CNIVX1 U4092 ( .A(n4102), .Z(n5144) );
  CNIVX1 U4093 ( .A(n5146), .Z(n5145) );
  CNIVX1 U4094 ( .A(n1565), .Z(n5146) );
  CNIVX1 U4095 ( .A(n5149), .Z(n5147) );
  CNIVX1 U4096 ( .A(n4115), .Z(n5148) );
  CENXL U4097 ( .A(opera2[57]), .B(n4479), .Z(n4116) );
  CNIVX1 U4098 ( .A(n1563), .Z(n5149) );
  CNIVX1 U4099 ( .A(n5152), .Z(n5150) );
  CNIVX1 U4100 ( .A(n4128), .Z(n5151) );
  CNIVX1 U4101 ( .A(n5153), .Z(n5152) );
  CNIVX1 U4102 ( .A(n1561), .Z(n5153) );
  CNIVX1 U4103 ( .A(n5156), .Z(n5154) );
  CNIVX1 U4104 ( .A(n4140), .Z(n5155) );
  CNIVX1 U4105 ( .A(n1559), .Z(n5156) );
  CEOXL U4106 ( .A(opera2[61]), .B(n4478), .Z(n4142) );
  CNR3XL U4107 ( .A(n5157), .B(n4148), .C(n4489), .Z(n3966) );
  CNR3XL U4108 ( .A(\cust[1] ), .B(n260), .C(n3479), .Z(n3483) );
  CNR3XL U4109 ( .A(n4148), .B(n1770), .C(n5157), .Z(n3949) );
  CIVX2 U4110 ( .A(n3775), .Z(n3165) );
  COND1XL U4111 ( .A(n3084), .B(n3104), .C(n3503), .Z(n3494) );
  COND1XL U4112 ( .A(n3094), .B(n3104), .C(n3503), .Z(n3550) );
  COND1XL U4113 ( .A(n3092), .B(n3104), .C(n3503), .Z(n3529) );
  COND1XL U4114 ( .A(n3090), .B(n3104), .C(n3503), .Z(n3509) );
  CND2X1 U4115 ( .A(n3124), .B(n3665), .Z(n3666) );
  CND2X1 U4116 ( .A(n3118), .B(n3687), .Z(n3688) );
  CND2X1 U4117 ( .A(n3112), .B(n3709), .Z(n3710) );
  CND3XL U4118 ( .A(n3134), .B(n3117), .C(n3692), .Z(n3693) );
  CND3XL U4119 ( .A(n3135), .B(n3111), .C(n3714), .Z(n3715) );
  CND3XL U4120 ( .A(n3132), .B(n3130), .C(n3654), .Z(n3655) );
  CND3XL U4121 ( .A(n3679), .B(n3120), .C(n3681), .Z(n3682) );
  CND3XL U4122 ( .A(n3701), .B(n3114), .C(n3703), .Z(n3704) );
  CND2X1 U4123 ( .A(n3122), .B(n3673), .Z(n3674) );
  CND2X1 U4124 ( .A(n3116), .B(n3695), .Z(n3696) );
  CND2X1 U4125 ( .A(n3110), .B(n3717), .Z(n3718) );
  CND2X1 U4126 ( .A(n3121), .B(n3676), .Z(n3677) );
  CND2X1 U4127 ( .A(n3115), .B(n3698), .Z(n3699) );
  CND2X1 U4128 ( .A(n3109), .B(n3720), .Z(n3721) );
  CND2X1 U4129 ( .A(n3108), .B(n3723), .Z(n3724) );
  CND2X1 U4130 ( .A(n3125), .B(n3662), .Z(n3663) );
  CND2X1 U4131 ( .A(n3119), .B(n3684), .Z(n3685) );
  CND2X1 U4132 ( .A(n3113), .B(n3706), .Z(n3707) );
  CND2X1 U4133 ( .A(n3107), .B(n3726), .Z(n3727) );
  COND1XL U4134 ( .A(n3098), .B(n3104), .C(n3503), .Z(n3590) );
  COND1XL U4135 ( .A(n3096), .B(n3104), .C(n3503), .Z(n3570) );
  CANR1XL U4136 ( .A(n3743), .B(n3744), .C(n3745), .Z(n3740) );
  CNR2X1 U4137 ( .A(n3082), .B(n3414), .Z(n3746) );
  CND3XL U4138 ( .A(n3173), .B(n3874), .C(n5181), .Z(n3879) );
  CND3XL U4139 ( .A(n3171), .B(n3895), .C(n3778), .Z(n3900) );
  CND3XL U4140 ( .A(n3175), .B(n3853), .C(n5182), .Z(n3858) );
  CND3XL U4141 ( .A(n3828), .B(n3832), .C(n3778), .Z(n3837) );
  CIVX2 U4142 ( .A(n3966), .Z(n3276) );
  CNR2X1 U4143 ( .A(n3738), .B(n3082), .Z(n3745) );
  CNR2X1 U4144 ( .A(n4480), .B(n4479), .Z(n3775) );
  COND1XL U4145 ( .A(n3126), .B(n3104), .C(n3503), .Z(n3630) );
  COND1XL U4146 ( .A(n3101), .B(n3104), .C(n3503), .Z(n3610) );
  CNIVX1 U4147 ( .A(n4168), .Z(n5186) );
  CNIVX1 U4148 ( .A(n4281), .Z(n5184) );
  CNR3XL U4149 ( .A(n3956), .B(n3964), .C(n3167), .Z(n3965) );
  CNR3XL U4150 ( .A(n3986), .B(n3992), .C(n3980), .Z(n3993) );
  CNR3XL U4151 ( .A(n4012), .B(n4018), .C(n4006), .Z(n4019) );
  CNR3XL U4152 ( .A(n4038), .B(n4044), .C(n4032), .Z(n4045) );
  CNR3XL U4153 ( .A(n4064), .B(n4070), .C(n4058), .Z(n4071) );
  CNR3XL U4154 ( .A(n4090), .B(n4096), .C(n4084), .Z(n4097) );
  CNR3XL U4155 ( .A(n4116), .B(n4122), .C(n4110), .Z(n4123) );
  CNR3XL U4156 ( .A(n3823), .B(n3827), .C(n3177), .Z(n3828) );
  CNR3XL U4157 ( .A(n3795), .B(n3799), .C(n3790), .Z(n3800) );
  CNR3XL U4158 ( .A(n3937), .B(n3946), .C(n3930), .Z(n3947) );
  CNR3XL U4159 ( .A(n3814), .B(n3818), .C(n3808), .Z(n3819) );
  CND3XL U4160 ( .A(n3972), .B(n3979), .C(n3965), .Z(n3980) );
  CND3XL U4161 ( .A(n3999), .B(n4005), .C(n3993), .Z(n4006) );
  CND3XL U4162 ( .A(n4025), .B(n4031), .C(n4019), .Z(n4032) );
  CND3XL U4163 ( .A(n4051), .B(n4057), .C(n4045), .Z(n4058) );
  CND3XL U4164 ( .A(n4077), .B(n4083), .C(n4071), .Z(n4084) );
  CND3XL U4165 ( .A(n4103), .B(n4109), .C(n4097), .Z(n4110) );
  CNR2X1 U4166 ( .A(n3774), .B(n3785), .Z(n3786) );
  CND3XL U4167 ( .A(n4129), .B(n4135), .C(n4123), .Z(n4136) );
  COND2X1 U4168 ( .A(\intadd_0/SUM[26] ), .B(n3278), .C(n4480), .D(n4687), .Z(
        n4132) );
  COND4CX1 U4169 ( .A(n4123), .B(n4129), .C(n4135), .D(n4136), .Z(n4134) );
  CANR2X1 U4170 ( .A(n4141), .B(n4481), .C(n5179), .D(n3209), .Z(n4140) );
  CANR1XL U4171 ( .A(n4142), .B(n4136), .C(n3765), .Z(n4141) );
  COND2X1 U4172 ( .A(n4485), .B(n3397), .C(\intadd_1/SUM[26] ), .D(n3277), .Z(
        n4130) );
  COND2X1 U4173 ( .A(n3391), .B(n4482), .C(\intadd_0/SUM[27] ), .D(n3275), .Z(
        n4131) );
  COND2X1 U4174 ( .A(\intadd_1/SUM[27] ), .B(n3276), .C(\intadd_1/SUM[28] ), 
        .D(n4487), .Z(n4133) );
  CANR2X1 U4175 ( .A(n4854), .B(n4481), .C(n3766), .D(n3233), .Z(n4068) );
  CANR4CX1 U4176 ( .A(n4064), .B(n4058), .C(n4070), .D(n4071), .Z(n4069) );
  CANR2X1 U4177 ( .A(n4807), .B(n4481), .C(n3766), .D(n3223), .Z(n4094) );
  CANR4CX1 U4178 ( .A(n4090), .B(n4084), .C(n4096), .D(n4097), .Z(n4095) );
  CANR2X1 U4179 ( .A(n4803), .B(n3647), .C(n3766), .D(n3213), .Z(n4120) );
  CANR4CX1 U4180 ( .A(n4116), .B(n4110), .C(n4122), .D(n4123), .Z(n4121) );
  CANR2X1 U4181 ( .A(n3647), .B(n5135), .C(n5179), .D(n3239), .Z(n4062) );
  CEOX1 U4182 ( .A(n4064), .B(n4058), .Z(n4063) );
  CANR2X1 U4183 ( .A(n4481), .B(n4076), .C(n5179), .D(n3234), .Z(n4075) );
  CEOX1 U4184 ( .A(n4071), .B(n4077), .Z(n4076) );
  CANR2X1 U4185 ( .A(n4481), .B(n4089), .C(n5179), .D(n3229), .Z(n4088) );
  CEOX1 U4186 ( .A(n4090), .B(n4084), .Z(n4089) );
  CANR2X1 U4187 ( .A(n4481), .B(n5144), .C(n5179), .D(n3224), .Z(n4101) );
  CEOX1 U4188 ( .A(n4097), .B(n4103), .Z(n4102) );
  CANR2X1 U4189 ( .A(n4481), .B(n5148), .C(n5179), .D(n3219), .Z(n4114) );
  CEOX1 U4190 ( .A(n4116), .B(n4110), .Z(n4115) );
  CANR2X1 U4191 ( .A(n3647), .B(n5151), .C(n5179), .D(n3214), .Z(n4127) );
  CEOX1 U4192 ( .A(n4123), .B(n4129), .Z(n4128) );
  CNR3XL U4193 ( .A(n5157), .B(n3206), .C(n4489), .Z(n3757) );
  COND2X1 U4194 ( .A(\intadd_0/SUM[14] ), .B(n3278), .C(n4480), .D(n4851), .Z(
        n4054) );
  COND4CX1 U4195 ( .A(n4045), .B(n4051), .C(n4057), .D(n4058), .Z(n4056) );
  COND2X1 U4196 ( .A(\intadd_0/SUM[18] ), .B(n3278), .C(n4480), .D(n4798), .Z(
        n4080) );
  COND4CX1 U4197 ( .A(n4071), .B(n4077), .C(n4083), .D(n4084), .Z(n4082) );
  COND2X1 U4198 ( .A(\intadd_0/SUM[22] ), .B(n3278), .C(n4480), .D(n4796), .Z(
        n4106) );
  COND4CX1 U4199 ( .A(n4097), .B(n4103), .C(n4109), .D(n4110), .Z(n4108) );
  COND2X1 U4200 ( .A(n4485), .B(n3236), .C(\intadd_1/SUM[14] ), .D(n3277), .Z(
        n4052) );
  COND2X1 U4201 ( .A(n3452), .B(n4482), .C(\intadd_0/SUM[15] ), .D(n3275), .Z(
        n4053) );
  COND2X1 U4202 ( .A(\intadd_1/SUM[15] ), .B(n3276), .C(\intadd_1/SUM[16] ), 
        .D(n4487), .Z(n4055) );
  COND2X1 U4203 ( .A(n4485), .B(n3226), .C(\intadd_1/SUM[18] ), .D(n3277), .Z(
        n4078) );
  COND2X1 U4204 ( .A(n3426), .B(n4482), .C(\intadd_0/SUM[19] ), .D(n3275), .Z(
        n4079) );
  COND2X1 U4205 ( .A(\intadd_1/SUM[19] ), .B(n3276), .C(\intadd_1/SUM[20] ), 
        .D(n4487), .Z(n4081) );
  COND2X1 U4206 ( .A(n4485), .B(n3216), .C(\intadd_1/SUM[22] ), .D(n3277), .Z(
        n4104) );
  COND2X1 U4207 ( .A(n3423), .B(n4482), .C(\intadd_0/SUM[23] ), .D(n3275), .Z(
        n4105) );
  COND2X1 U4208 ( .A(\intadd_1/SUM[23] ), .B(n3276), .C(\intadd_1/SUM[24] ), 
        .D(n4487), .Z(n4107) );
  CNR2X1 U4209 ( .A(n3138), .B(n3497), .Z(n3489) );
  CANR2X1 U4210 ( .A(n4858), .B(n3647), .C(n3766), .D(n3243), .Z(n4042) );
  CANR4CX1 U4211 ( .A(n4038), .B(n4032), .C(n4044), .D(n4045), .Z(n4043) );
  CANR2X1 U4212 ( .A(n4963), .B(n3647), .C(n3766), .D(n3263), .Z(n3990) );
  CANR4CX1 U4213 ( .A(n3986), .B(n3980), .C(n3992), .D(n3993), .Z(n3991) );
  CANR2X1 U4214 ( .A(n4915), .B(n3647), .C(n3766), .D(n3253), .Z(n4016) );
  CANR4CX1 U4215 ( .A(n4012), .B(n4006), .C(n4018), .D(n4019), .Z(n4017) );
  CANR2X1 U4216 ( .A(n3647), .B(n5116), .C(n5179), .D(n3269), .Z(n3984) );
  CEOX1 U4217 ( .A(n3986), .B(n3980), .Z(n3985) );
  CANR2X1 U4218 ( .A(n3647), .B(n3998), .C(n5179), .D(n3264), .Z(n3997) );
  CEOX1 U4219 ( .A(n3993), .B(n3999), .Z(n3998) );
  CANR2X1 U4220 ( .A(n3647), .B(n5122), .C(n5179), .D(n3259), .Z(n4010) );
  CEOX1 U4221 ( .A(n4012), .B(n4006), .Z(n4011) );
  CANR2X1 U4222 ( .A(n3647), .B(n5125), .C(n5179), .D(n3254), .Z(n4023) );
  CEOX1 U4223 ( .A(n4019), .B(n4025), .Z(n4024) );
  CANR2X1 U4224 ( .A(n3647), .B(n5129), .C(n5179), .D(n3249), .Z(n4036) );
  CEOX1 U4225 ( .A(n4038), .B(n4032), .Z(n4037) );
  CANR2X1 U4226 ( .A(n3647), .B(n4050), .C(n5179), .D(n3244), .Z(n4049) );
  CEOX1 U4227 ( .A(n4045), .B(n4051), .Z(n4050) );
  COND2X1 U4228 ( .A(\intadd_0/SUM[6] ), .B(n3278), .C(n4480), .D(n4912), .Z(
        n4002) );
  COND4CX1 U4229 ( .A(n3993), .B(n3999), .C(n4005), .D(n4006), .Z(n4004) );
  COND2X1 U4230 ( .A(\intadd_0/SUM[10] ), .B(n3278), .C(n4480), .D(n4910), .Z(
        n4028) );
  COND4CX1 U4231 ( .A(n4019), .B(n4025), .C(n4031), .D(n4032), .Z(n4030) );
  COND2X1 U4232 ( .A(\intadd_0/SUM[2] ), .B(n3278), .C(n4480), .D(n4994), .Z(
        n3976) );
  COND4CX1 U4233 ( .A(n3965), .B(n3972), .C(n3979), .D(n3980), .Z(n3978) );
  COND2X1 U4234 ( .A(\intadd_1/SUM[7] ), .B(n3276), .C(\intadd_1/SUM[8] ), .D(
        n4487), .Z(n4003) );
  COND2X1 U4235 ( .A(n4485), .B(n3256), .C(\intadd_1/SUM[6] ), .D(n3277), .Z(
        n4000) );
  COND2X1 U4236 ( .A(n3466), .B(n4482), .C(\intadd_0/SUM[7] ), .D(n3275), .Z(
        n4001) );
  COND2X1 U4237 ( .A(n4485), .B(n3246), .C(\intadd_1/SUM[10] ), .D(n3277), .Z(
        n4026) );
  COND2X1 U4238 ( .A(n3464), .B(n4482), .C(\intadd_0/SUM[11] ), .D(n3275), .Z(
        n4027) );
  COND2X1 U4239 ( .A(\intadd_1/SUM[11] ), .B(n3276), .C(\intadd_1/SUM[12] ), 
        .D(n4487), .Z(n4029) );
  CENX1 U4240 ( .A(n3136), .B(n3162), .Z(n3657) );
  CENX1 U4241 ( .A(n3136), .B(n3163), .Z(n3654) );
  CENX1 U4242 ( .A(n3136), .B(n4919), .Z(n3673) );
  CENX1 U4243 ( .A(n3136), .B(n4967), .Z(n3662) );
  CENX1 U4244 ( .A(n3136), .B(n3160), .Z(n3665) );
  COND1XL U4245 ( .A(n3533), .B(n3200), .C(n3545), .Z(n3539) );
  CANR4CX1 U4246 ( .A(n4486), .B(n3533), .C(n3539), .D(n4815), .Z(n3538) );
  CANR4CX1 U4247 ( .A(n3937), .B(n3930), .C(n3946), .D(n3947), .Z(n3941) );
  CANR2X1 U4248 ( .A(n4959), .B(n4481), .C(n3766), .D(n3313), .Z(n3962) );
  CANR4CX1 U4249 ( .A(n3956), .B(n3167), .C(n3964), .D(n3965), .Z(n3963) );
  CANR2X1 U4250 ( .A(n3647), .B(n3954), .C(n5179), .D(n3476), .Z(n3953) );
  CENX1 U4251 ( .A(n3956), .B(n3947), .Z(n3954) );
  CANR2X1 U4252 ( .A(n3647), .B(n5113), .C(n5179), .D(n3314), .Z(n3970) );
  CEOX1 U4253 ( .A(n3965), .B(n3972), .Z(n3971) );
  COND2X1 U4254 ( .A(n3401), .B(n4481), .C(n4480), .D(n3713), .Z(n1662) );
  COND4CX1 U4255 ( .A(n3111), .B(n3135), .C(n3714), .D(n3715), .Z(n3713) );
  COND2X1 U4256 ( .A(n3385), .B(n4481), .C(n4480), .D(n3731), .Z(n1656) );
  CENX1 U4257 ( .A(n3730), .B(n3732), .Z(n3731) );
  CND3XL U4258 ( .A(n3133), .B(n3123), .C(n3670), .Z(n3671) );
  CND3XL U4259 ( .A(n3657), .B(n3129), .C(n3659), .Z(n3660) );
  COND4CX1 U4260 ( .A(n5192), .B(n3533), .C(n3537), .D(n4815), .Z(n3536) );
  CNR2X1 U4261 ( .A(n3533), .B(n3103), .Z(n3537) );
  CEOX1 U4262 ( .A(n3930), .B(n3937), .Z(n3936) );
  COND1XL U4263 ( .A(n3400), .B(n4481), .C(n3708), .Z(n1664) );
  COND3X1 U4264 ( .A(n3112), .B(n3709), .C(n3710), .D(n3647), .Z(n3708) );
  COND1XL U4265 ( .A(n3384), .B(n3647), .C(n3725), .Z(n1658) );
  COND3X1 U4266 ( .A(n3107), .B(n3726), .C(n3727), .D(n4481), .Z(n3725) );
  COND1XL U4267 ( .A(n3383), .B(n3647), .C(n3719), .Z(n1660) );
  COND3X1 U4268 ( .A(n3109), .B(n3720), .C(n3721), .D(n3647), .Z(n3719) );
  CND4X1 U4269 ( .A(n3968), .B(n3271), .C(n3969), .D(n3970), .Z(n1585) );
  CANR2X1 U4270 ( .A(n5187), .B(n3268), .C(n4484), .D(n3270), .Z(n3968) );
  CANR2X1 U4271 ( .A(n5178), .B(n3312), .C(n5190), .D(n3269), .Z(n3969) );
  CNR3XL U4272 ( .A(n5157), .B(n3944), .C(n4489), .Z(n3967) );
  CNR2X1 U4273 ( .A(n3752), .B(n3082), .Z(n3738) );
  CND2X1 U4274 ( .A(n4174), .B(n3439), .Z(n3944) );
  CENX1 U4275 ( .A(n3136), .B(n3156), .Z(n3679) );
  CNR3XL U4276 ( .A(n4165), .B(n3483), .C(n4166), .Z(n3753) );
  CENX1 U4277 ( .A(n3136), .B(n3151), .Z(n3692) );
  CENX1 U4278 ( .A(n3136), .B(n3155), .Z(n3681) );
  CANR1XL U4279 ( .A(n3361), .B(n3414), .C(n3082), .Z(n3735) );
  CENX1 U4280 ( .A(n3136), .B(n4866), .Z(n3695) );
  CENX1 U4281 ( .A(n3136), .B(n3157), .Z(n3676) );
  CENX1 U4282 ( .A(n3136), .B(n3149), .Z(n3698) );
  CENX1 U4283 ( .A(n3136), .B(n4862), .Z(n3684) );
  CENX1 U4284 ( .A(n3136), .B(n3153), .Z(n3687) );
  CNR2X1 U4285 ( .A(n4150), .B(n3944), .Z(n4165) );
  COND1XL U4286 ( .A(n3576), .B(n3200), .C(n3545), .Z(n3580) );
  COND1XL U4287 ( .A(n3556), .B(n3200), .C(n3545), .Z(n3560) );
  CANR4CX1 U4288 ( .A(n4486), .B(n3576), .C(n3580), .D(n4862), .Z(n3579) );
  CANR4CX1 U4289 ( .A(n4486), .B(n3556), .C(n3560), .D(n4866), .Z(n3559) );
  COND2X1 U4290 ( .A(n3945), .B(n3276), .C(\intadd_1/SUM[0] ), .D(n4487), .Z(
        n3942) );
  CAN8X1 U4291 ( .A(n3433), .B(n3422), .C(n3421), .D(n3409), .E(n3434), .F(
        n3431), .G(n4276), .H(n4277), .Z(n4174) );
  CAN6X1 U4292 ( .A(n3428), .B(n3416), .C(n3412), .D(n3417), .E(n3435), .F(
        n3436), .Z(n4276) );
  CAN8X1 U4293 ( .A(n3411), .B(n3427), .C(n3410), .D(n3429), .E(n3425), .F(
        n3407), .G(n3418), .H(n4278), .Z(n4277) );
  CAN6X1 U4294 ( .A(n3432), .B(n3419), .C(n3408), .D(n3420), .E(n3395), .F(
        n3430), .Z(n4278) );
  COND2X1 U4295 ( .A(n3459), .B(n4481), .C(n4480), .D(n3680), .Z(n1674) );
  COND4CX1 U4296 ( .A(n3120), .B(n3679), .C(n3681), .D(n3682), .Z(n3680) );
  COND2X1 U4297 ( .A(n3444), .B(n4481), .C(n4480), .D(n3691), .Z(n1670) );
  COND2X1 U4298 ( .A(n3399), .B(n4481), .C(n4480), .D(n3702), .Z(n1666) );
  COND4CX1 U4299 ( .A(n3114), .B(n3701), .C(n3703), .D(n3704), .Z(n3702) );
  CND3XL U4300 ( .A(n3172), .B(n3884), .C(n3778), .Z(n3889) );
  CND3XL U4301 ( .A(n3174), .B(n3863), .C(n5181), .Z(n3868) );
  CND3XL U4302 ( .A(n3176), .B(n3842), .C(n5182), .Z(n3847) );
  CND2X1 U4303 ( .A(n3751), .B(n3743), .Z(n3749) );
  COND4CX1 U4304 ( .A(n5192), .B(n3576), .C(n3578), .D(n4862), .Z(n3577) );
  CNR2X1 U4305 ( .A(n3576), .B(n3103), .Z(n3578) );
  COND4CX1 U4306 ( .A(n5192), .B(n3556), .C(n3558), .D(n4866), .Z(n3557) );
  CNR2X1 U4307 ( .A(n3556), .B(n3103), .Z(n3558) );
  CNR2X1 U4308 ( .A(n3772), .B(n3291), .Z(n3771) );
  CNR2X1 U4309 ( .A(n4150), .B(n4148), .Z(n4177) );
  COND1XL U4310 ( .A(n3445), .B(n4481), .C(n3697), .Z(n1668) );
  COND3X1 U4311 ( .A(n3115), .B(n3698), .C(n3699), .D(n4481), .Z(n3697) );
  COND1XL U4312 ( .A(n3443), .B(n4481), .C(n3686), .Z(n1672) );
  COND3X1 U4313 ( .A(n3118), .B(n3687), .C(n3688), .D(n4481), .Z(n3686) );
  COND1XL U4314 ( .A(n3743), .B(n3361), .C(n3747), .Z(n1625) );
  CANR1XL U4315 ( .A(n3738), .B(n3361), .C(n3083), .Z(n3747) );
  COR2X1 U4316 ( .A(n3758), .B(n5191), .Z(n5157) );
  CNR2X1 U4317 ( .A(n3745), .B(n3436), .Z(n1637) );
  CNR2X1 U4318 ( .A(n3743), .B(n3435), .Z(n1635) );
  CNR2X1 U4319 ( .A(n3745), .B(n3434), .Z(n1641) );
  CNR2X1 U4320 ( .A(n3745), .B(n3433), .Z(n1645) );
  CNR2X1 U4321 ( .A(n3745), .B(n3432), .Z(n1633) );
  CNR2X1 U4322 ( .A(n3743), .B(n3431), .Z(n1643) );
  CNR2X1 U4323 ( .A(n3743), .B(n3430), .Z(n1631) );
  CNR2X1 U4324 ( .A(n3743), .B(n3429), .Z(n1647) );
  CNR2X1 U4325 ( .A(n3743), .B(n3428), .Z(n1639) );
  CNR2X1 U4326 ( .A(n3745), .B(n3427), .Z(n1649) );
  CNR2X1 U4327 ( .A(n3745), .B(n3425), .Z(n1627) );
  CNR2X1 U4328 ( .A(n3745), .B(n3422), .Z(n1644) );
  CNR2X1 U4329 ( .A(n3743), .B(n3421), .Z(n1646) );
  CNR2X1 U4330 ( .A(n3743), .B(n3420), .Z(n1630) );
  CNR2X1 U4331 ( .A(n3745), .B(n3419), .Z(n1632) );
  CNR2X1 U4332 ( .A(n3745), .B(n3418), .Z(n1628) );
  CNR2X1 U4333 ( .A(n3745), .B(n3417), .Z(n1636) );
  CNR2X1 U4334 ( .A(n3743), .B(n3416), .Z(n1638) );
  CNR2X1 U4335 ( .A(n3745), .B(n3412), .Z(n1640) );
  CNR2X1 U4336 ( .A(n3746), .B(n3411), .Z(n1650) );
  CNR2X1 U4337 ( .A(n3745), .B(n3410), .Z(n1648) );
  CNR2X1 U4338 ( .A(n3743), .B(n3409), .Z(n1642) );
  CNR2X1 U4339 ( .A(n3743), .B(n3408), .Z(n1634) );
  CNR2X1 U4340 ( .A(n3745), .B(n3407), .Z(n1626) );
  CNR2X1 U4341 ( .A(n3745), .B(n3395), .Z(n1629) );
  CND2X1 U4342 ( .A(n5191), .B(n3754), .Z(n3743) );
  CANR1XL U4343 ( .A(n3136), .B(n3200), .C(n4476), .Z(n3492) );
  CENX1 U4344 ( .A(n3136), .B(n3148), .Z(n3701) );
  CNR3XL U4345 ( .A(n3078), .B(n3475), .C(n4170), .Z(n4309) );
  CNR2X1 U4346 ( .A(n4476), .B(n4478), .Z(n3777) );
  CNR2X1 U4347 ( .A(n3200), .B(n4476), .Z(n3647) );
  CND3XL U4348 ( .A(n4468), .B(n3475), .C(n3415), .Z(n4281) );
  CENX1 U4349 ( .A(n3136), .B(n3143), .Z(n3714) );
  CENX1 U4350 ( .A(n3136), .B(n3147), .Z(n3703) );
  CENX1 U4351 ( .A(n3136), .B(n3142), .Z(n3717) );
  CENX1 U4352 ( .A(n3136), .B(n3141), .Z(n3720) );
  CENX1 U4353 ( .A(n3136), .B(n3140), .Z(n3723) );
  CENX1 U4354 ( .A(n3136), .B(n4815), .Z(n3706) );
  CENX1 U4355 ( .A(n3136), .B(n3139), .Z(n3726) );
  CENX1 U4356 ( .A(n3136), .B(n3145), .Z(n3709) );
  CENX1 U4357 ( .A(n4479), .B(n3194), .Z(n3832) );
  CENX1 U4358 ( .A(n4479), .B(n3191), .Z(n3853) );
  CENX1 U4359 ( .A(n4479), .B(n3185), .Z(n3895) );
  CENX1 U4360 ( .A(n4479), .B(n3188), .Z(n3874) );
  CIVX2 U4361 ( .A(n3488), .Z(n3103) );
  CENX1 U4362 ( .A(n4479), .B(n3182), .Z(n3916) );
  COND1XL U4363 ( .A(n3616), .B(n3200), .C(n3545), .Z(n3620) );
  COND1XL U4364 ( .A(n3596), .B(n3200), .C(n3545), .Z(n3600) );
  CANR4CX1 U4365 ( .A(n4486), .B(n3596), .C(n3600), .D(n4919), .Z(n3599) );
  COND1XL U4366 ( .A(n3635), .B(n3104), .C(n3503), .Z(n3640) );
  CNR3XL U4367 ( .A(n3440), .B(n3361), .C(n3437), .Z(n3744) );
  CANR1XL U4368 ( .A(n4478), .B(n3200), .C(n4476), .Z(n5182) );
  CANR1XL U4369 ( .A(n4478), .B(n3200), .C(n4476), .Z(n5181) );
  CANR1XL U4370 ( .A(n4478), .B(n3200), .C(n4476), .Z(n3778) );
  CND2X1 U4371 ( .A(n3545), .B(n3200), .Z(n3503) );
  COND1XL U4372 ( .A(n4170), .B(n3389), .C(n3754), .Z(n4468) );
  CND2X1 U4373 ( .A(n4179), .B(n4489), .Z(n4143) );
  COND2X1 U4374 ( .A(n3469), .B(n4481), .C(n4480), .D(n3658), .Z(n1682) );
  COND2X1 U4375 ( .A(n3468), .B(n4481), .C(n4480), .D(n3653), .Z(n1684) );
  COND4CX1 U4376 ( .A(n3130), .B(n3132), .C(n3654), .D(n3655), .Z(n3653) );
  COND2X1 U4377 ( .A(n3457), .B(n4481), .C(n4480), .D(n3669), .Z(n1678) );
  COND4CX1 U4378 ( .A(n3123), .B(n3133), .C(n3670), .D(n3671), .Z(n3669) );
  CNR2X1 U4379 ( .A(n3616), .B(n3103), .Z(n3618) );
  CIVX2 U4380 ( .A(n3545), .Z(n3104) );
  CNR2X1 U4381 ( .A(n3758), .B(n4148), .Z(n4179) );
  CND3XL U4382 ( .A(n3800), .B(n3804), .C(n3778), .Z(n3809) );
  COND4CX1 U4383 ( .A(n5192), .B(n3616), .C(n3618), .D(n4967), .Z(n3617) );
  CANR4CX1 U4384 ( .A(n4486), .B(n3616), .C(n3620), .D(n4967), .Z(n3619) );
  COND4CX1 U4385 ( .A(n5192), .B(n3596), .C(n3598), .D(n4919), .Z(n3597) );
  CNR2X1 U4386 ( .A(n3596), .B(n3103), .Z(n3598) );
  COND1XL U4387 ( .A(n3475), .B(n4477), .C(n3645), .Z(n224) );
  CANR2X1 U4388 ( .A(n3545), .B(n4479), .C(n5192), .D(n4478), .Z(n3645) );
  COND1XL U4389 ( .A(n3458), .B(n4481), .C(n3675), .Z(n1676) );
  COND3X1 U4390 ( .A(n3121), .B(n3676), .C(n3677), .D(n4481), .Z(n3675) );
  COND1XL U4391 ( .A(n3456), .B(n4481), .C(n3664), .Z(n1680) );
  COND3X1 U4392 ( .A(n3124), .B(n3665), .C(n3666), .D(n3647), .Z(n3664) );
  CND2X1 U4393 ( .A(n3777), .B(n3195), .Z(n3810) );
  CND2X1 U4394 ( .A(n3777), .B(n3186), .Z(n3890) );
  CND2X1 U4395 ( .A(n3777), .B(n3187), .Z(n3880) );
  CND2X1 U4396 ( .A(n3777), .B(n3189), .Z(n3869) );
  CND2X1 U4397 ( .A(n3777), .B(n3192), .Z(n3848) );
  CND2X1 U4398 ( .A(n3777), .B(n3184), .Z(n3901) );
  CND2X1 U4399 ( .A(n3777), .B(n3190), .Z(n3859) );
  CND2X1 U4400 ( .A(n3777), .B(n3193), .Z(n3838) );
  CAN2X1 U4401 ( .A(n3767), .B(n4481), .Z(n3764) );
  CENX1 U4402 ( .A(n3136), .B(n3138), .Z(n3729) );
  COND3X1 U4403 ( .A(n3392), .B(n4281), .C(n4451), .D(n4452), .Z(n1432) );
  CND2X1 U4404 ( .A(result[58]), .B(n3078), .Z(n4452) );
  COND3X1 U4405 ( .A(result_not[58]), .B(n3301), .C(n4453), .D(n4475), .Z(
        n4451) );
  COND3X1 U4406 ( .A(n3221), .B(n5184), .C(n4442), .D(n4443), .Z(n1435) );
  CND2X1 U4407 ( .A(result[55]), .B(n3078), .Z(n4443) );
  COND3X1 U4408 ( .A(n3304), .B(result_not[55]), .C(n4444), .D(n5183), .Z(
        n4442) );
  CND3XL U4409 ( .A(result_not[1]), .B(result_not[0]), .C(cina), .Z(n4285) );
  CND3XL U4410 ( .A(result_not[3]), .B(result_not[2]), .C(n3359), .Z(n4290) );
  CND3XL U4411 ( .A(result_not[5]), .B(result_not[4]), .C(n3358), .Z(n4295) );
  CND3XL U4412 ( .A(result_not[7]), .B(result_not[6]), .C(n3357), .Z(n4300) );
  CND3XL U4413 ( .A(result_not[9]), .B(result_not[8]), .C(n3356), .Z(n4305) );
  CND2X1 U4414 ( .A(n3292), .B(result_not[62]), .Z(n4465) );
  COND3X1 U4415 ( .A(n3393), .B(n4281), .C(n4463), .D(n4464), .Z(n1428) );
  CND2X1 U4416 ( .A(result[62]), .B(n3078), .Z(n4464) );
  COND3X1 U4417 ( .A(result_not[62]), .B(n3292), .C(n4465), .D(n4475), .Z(
        n4463) );
  COND3X1 U4418 ( .A(n3391), .B(n4281), .C(n4457), .D(n4458), .Z(n1430) );
  CND2X1 U4419 ( .A(result[60]), .B(n3078), .Z(n4458) );
  COND3X1 U4420 ( .A(result_not[60]), .B(n3299), .C(n4459), .D(n5183), .Z(
        n4457) );
  COND3X1 U4421 ( .A(n3423), .B(n5184), .C(n4445), .D(n4446), .Z(n1434) );
  CND2X1 U4422 ( .A(result[56]), .B(n3078), .Z(n4446) );
  COND3X1 U4423 ( .A(result_not[56]), .B(n3303), .C(n4447), .D(n5183), .Z(
        n4445) );
  COND3X1 U4424 ( .A(n3397), .B(n4281), .C(n4460), .D(n4461), .Z(n1429) );
  CND2X1 U4425 ( .A(result[61]), .B(n3078), .Z(n4461) );
  COND3X1 U4426 ( .A(n3298), .B(result_not[61]), .C(n4462), .D(n5183), .Z(
        n4460) );
  COND3X1 U4427 ( .A(n3211), .B(n4281), .C(n4454), .D(n4455), .Z(n1431) );
  CND2X1 U4428 ( .A(result[59]), .B(n3078), .Z(n4455) );
  COND3X1 U4429 ( .A(n3300), .B(result_not[59]), .C(n4456), .D(n5183), .Z(
        n4454) );
  COND3X1 U4430 ( .A(n3216), .B(n5184), .C(n4448), .D(n4449), .Z(n1433) );
  CND2X1 U4431 ( .A(result[57]), .B(n3078), .Z(n4449) );
  COND3X1 U4432 ( .A(n3302), .B(result_not[57]), .C(n4450), .D(n4475), .Z(
        n4448) );
  CND2X1 U4433 ( .A(n3355), .B(result_not[10]), .Z(n4308) );
  CND2X1 U4434 ( .A(n3354), .B(result_not[11]), .Z(n4312) );
  CND2X1 U4435 ( .A(n3353), .B(result_not[12]), .Z(n4315) );
  CND2X1 U4436 ( .A(n3352), .B(result_not[13]), .Z(n4318) );
  CND2X1 U4437 ( .A(n3351), .B(result_not[14]), .Z(n4321) );
  CND2X1 U4438 ( .A(n3350), .B(result_not[15]), .Z(n4324) );
  CND2X1 U4439 ( .A(n3349), .B(result_not[16]), .Z(n4327) );
  CND2X1 U4440 ( .A(n3348), .B(result_not[17]), .Z(n4330) );
  CND2X1 U4441 ( .A(n3347), .B(result_not[18]), .Z(n4333) );
  CND2X1 U4442 ( .A(n3346), .B(result_not[19]), .Z(n4336) );
  CND2X1 U4443 ( .A(n3345), .B(result_not[20]), .Z(n4339) );
  CND2X1 U4444 ( .A(n3344), .B(result_not[21]), .Z(n4342) );
  CND2X1 U4445 ( .A(n3343), .B(result_not[22]), .Z(n4345) );
  CND2X1 U4446 ( .A(n3342), .B(result_not[23]), .Z(n4348) );
  CND2X1 U4447 ( .A(n3341), .B(result_not[24]), .Z(n4351) );
  CND2X1 U4448 ( .A(n3340), .B(result_not[25]), .Z(n4354) );
  CND2X1 U4449 ( .A(n3339), .B(result_not[26]), .Z(n4357) );
  CND2X1 U4450 ( .A(n3338), .B(result_not[27]), .Z(n4360) );
  CND2X1 U4451 ( .A(n3337), .B(result_not[28]), .Z(n4363) );
  CND2X1 U4452 ( .A(n3336), .B(result_not[29]), .Z(n4366) );
  CND2X1 U4453 ( .A(n3335), .B(result_not[30]), .Z(n4369) );
  CND2X1 U4454 ( .A(n3334), .B(result_not[31]), .Z(n4372) );
  CND2X1 U4455 ( .A(n3333), .B(result_not[32]), .Z(n4375) );
  CND2X1 U4456 ( .A(n3332), .B(result_not[33]), .Z(n4378) );
  CND2X1 U4457 ( .A(n3331), .B(result_not[34]), .Z(n4381) );
  CND2X1 U4458 ( .A(n3330), .B(result_not[35]), .Z(n4384) );
  CND2X1 U4459 ( .A(n3329), .B(result_not[36]), .Z(n4387) );
  CND2X1 U4460 ( .A(n3328), .B(result_not[37]), .Z(n4390) );
  CND2X1 U4461 ( .A(n3327), .B(result_not[38]), .Z(n4393) );
  CND2X1 U4462 ( .A(n3326), .B(result_not[39]), .Z(n4396) );
  CND2X1 U4463 ( .A(n3325), .B(result_not[40]), .Z(n4399) );
  CND2X1 U4464 ( .A(n3324), .B(result_not[41]), .Z(n4402) );
  CND2X1 U4465 ( .A(n3323), .B(result_not[42]), .Z(n4405) );
  CND2X1 U4466 ( .A(n3322), .B(result_not[43]), .Z(n4408) );
  CND2X1 U4467 ( .A(n3321), .B(result_not[44]), .Z(n4411) );
  CND2X1 U4468 ( .A(n3320), .B(result_not[45]), .Z(n4414) );
  CND2X1 U4469 ( .A(n3319), .B(result_not[46]), .Z(n4417) );
  CND2X1 U4470 ( .A(n3318), .B(result_not[47]), .Z(n4420) );
  CND2X1 U4471 ( .A(n3311), .B(result_not[48]), .Z(n4423) );
  CND2X1 U4472 ( .A(n3310), .B(result_not[49]), .Z(n4426) );
  CND2X1 U4473 ( .A(n3309), .B(result_not[50]), .Z(n4429) );
  CND2X1 U4474 ( .A(n3308), .B(result_not[51]), .Z(n4432) );
  CND2X1 U4475 ( .A(n3307), .B(result_not[52]), .Z(n4435) );
  CND2X1 U4476 ( .A(n3306), .B(result_not[53]), .Z(n4438) );
  CND2X1 U4477 ( .A(n3305), .B(result_not[54]), .Z(n4441) );
  CND2X1 U4478 ( .A(n3304), .B(result_not[55]), .Z(n4444) );
  CND2X1 U4479 ( .A(n3303), .B(result_not[56]), .Z(n4447) );
  CND2X1 U4480 ( .A(n3302), .B(result_not[57]), .Z(n4450) );
  CND2X1 U4481 ( .A(n3301), .B(result_not[58]), .Z(n4453) );
  CND2X1 U4482 ( .A(n3300), .B(result_not[59]), .Z(n4456) );
  CND2X1 U4483 ( .A(n3299), .B(result_not[60]), .Z(n4459) );
  CND2X1 U4484 ( .A(n3298), .B(result_not[61]), .Z(n4462) );
  COND2X1 U4485 ( .A(n3396), .B(n4281), .C(n4467), .D(n4474), .Z(n4466) );
  CEOX1 U4486 ( .A(n4465), .B(result_not[63]), .Z(n4467) );
  CND2X1 U4487 ( .A(n4161), .B(n3800), .Z(n3808) );
  CANR4CX1 U4488 ( .A(n4479), .B(n3196), .C(n4521), .D(n4163), .Z(n4161) );
  CANR1XL U4489 ( .A(n4479), .B(n3196), .C(n4521), .Z(n4163) );
  CND2X1 U4490 ( .A(n4151), .B(n3168), .Z(n3930) );
  CANR4CX1 U4491 ( .A(n4479), .B(n3181), .C(n4528), .D(n4164), .Z(n4151) );
  CANR1XL U4492 ( .A(n4479), .B(n3181), .C(n4528), .Z(n4164) );
  CENX1 U4493 ( .A(n4478), .B(n4524), .Z(n4162) );
  CENX1 U4494 ( .A(n4479), .B(n5046), .Z(n3785) );
  COND3X1 U4495 ( .A(n4517), .B(n3891), .C(n4155), .D(n3172), .Z(n3888) );
  COND3X1 U4496 ( .A(n4513), .B(n3870), .C(n4157), .D(n3174), .Z(n3867) );
  COND3X1 U4497 ( .A(n4511), .B(n3849), .C(n4159), .D(n3176), .Z(n3846) );
  COND3X1 U4498 ( .A(n4501), .B(n3912), .C(n4153), .D(n3170), .Z(n3909) );
  COND1XL U4499 ( .A(n4479), .B(n3183), .C(n4501), .Z(n4153) );
  COND3X1 U4500 ( .A(n4479), .B(n4519), .C(n3169), .D(n4152), .Z(n3920) );
  CANR2X1 U4501 ( .A(n4519), .B(n3182), .C(n5090), .D(n4479), .Z(n4152) );
  COND3X1 U4502 ( .A(n4479), .B(n4515), .C(n3173), .D(n4156), .Z(n3878) );
  CANR2X1 U4503 ( .A(n4515), .B(n3188), .C(n5068), .D(n4479), .Z(n4156) );
  COND3X1 U4504 ( .A(n4479), .B(n4507), .C(n3171), .D(n4154), .Z(n3899) );
  CANR2X1 U4505 ( .A(n4507), .B(n3185), .C(n5079), .D(n4479), .Z(n4154) );
  COND3X1 U4506 ( .A(n4479), .B(n4505), .C(n3175), .D(n4158), .Z(n3857) );
  CANR2X1 U4507 ( .A(n4505), .B(n3191), .C(n5058), .D(n4479), .Z(n4158) );
  COND3X1 U4508 ( .A(n4479), .B(n4503), .C(n3828), .D(n4160), .Z(n3836) );
  CANR2X1 U4509 ( .A(n4503), .B(n3194), .C(n4539), .D(n4479), .Z(n4160) );
  CANR2X1 U4510 ( .A(n4481), .B(n4149), .C(n5188), .D(D[31]), .Z(n4145) );
  CEOX1 U4511 ( .A(n3765), .B(n3767), .Z(n4149) );
  CND2X1 U4512 ( .A(cin2a), .B(n3780), .Z(n3774) );
  CANR1XL U4513 ( .A(D[31]), .B(n4483), .C(n3762), .Z(n3761) );
  CANR2X1 U4514 ( .A(n3764), .B(n3765), .C(n3766), .D(n3202), .Z(n3760) );
  COND2X1 U4515 ( .A(n3763), .B(n3275), .C(\intadd_1/SUM[29] ), .D(n3277), .Z(
        n3762) );
  COND3X1 U4516 ( .A(n3424), .B(n5184), .C(n4439), .D(n4440), .Z(n1436) );
  CND2X1 U4517 ( .A(result[54]), .B(n3078), .Z(n4440) );
  COND3X1 U4518 ( .A(result_not[54]), .B(n3305), .C(n4441), .D(n4309), .Z(
        n4439) );
  COND3X1 U4519 ( .A(n3426), .B(n5184), .C(n4433), .D(n4434), .Z(n1438) );
  CND2X1 U4520 ( .A(result[52]), .B(n3078), .Z(n4434) );
  COND3X1 U4521 ( .A(result_not[52]), .B(n3307), .C(n4435), .D(n4475), .Z(
        n4433) );
  COND3X1 U4522 ( .A(n3451), .B(n5184), .C(n4427), .D(n4428), .Z(n1440) );
  CND2X1 U4523 ( .A(result[50]), .B(n3078), .Z(n4428) );
  COND3X1 U4524 ( .A(result_not[50]), .B(n3309), .C(n4429), .D(n5183), .Z(
        n4427) );
  COND3X1 U4525 ( .A(n3452), .B(n5184), .C(n4421), .D(n4422), .Z(n1442) );
  CND2X1 U4526 ( .A(result[48]), .B(n3078), .Z(n4422) );
  COND3X1 U4527 ( .A(result_not[48]), .B(n3311), .C(n4423), .D(n4309), .Z(
        n4421) );
  COND3X1 U4528 ( .A(n3226), .B(n5184), .C(n4436), .D(n4437), .Z(n1437) );
  CND2X1 U4529 ( .A(result[53]), .B(n3078), .Z(n4437) );
  COND3X1 U4530 ( .A(n3306), .B(result_not[53]), .C(n4438), .D(n4475), .Z(
        n4436) );
  COND3X1 U4531 ( .A(n3231), .B(n5184), .C(n4430), .D(n4431), .Z(n1439) );
  CND2X1 U4532 ( .A(result[51]), .B(n3078), .Z(n4431) );
  COND3X1 U4533 ( .A(n3308), .B(result_not[51]), .C(n4432), .D(n4475), .Z(
        n4430) );
  COND3X1 U4534 ( .A(n3236), .B(n5184), .C(n4424), .D(n4425), .Z(n1441) );
  CND2X1 U4535 ( .A(result[49]), .B(n3078), .Z(n4425) );
  COND3X1 U4536 ( .A(n3310), .B(result_not[49]), .C(n4426), .D(n4309), .Z(
        n4424) );
  COND3X1 U4537 ( .A(n3241), .B(n5184), .C(n4418), .D(n4419), .Z(n1443) );
  CND2X1 U4538 ( .A(result[47]), .B(n3078), .Z(n4419) );
  COND3X1 U4539 ( .A(n3318), .B(result_not[47]), .C(n4420), .D(n4475), .Z(
        n4418) );
  CANR2X1 U4540 ( .A(n5188), .B(D[30]), .C(n1734), .D(n5191), .Z(n4138) );
  CANR2X1 U4541 ( .A(n5187), .B(n3203), .C(n4484), .D(n3208), .Z(n4137) );
  CANR2X1 U4542 ( .A(n5178), .B(n3204), .C(n5190), .D(n3207), .Z(n4139) );
  CANR2X1 U4543 ( .A(n3949), .B(n3202), .C(n4483), .D(D[30]), .Z(n4144) );
  CANR2X1 U4544 ( .A(n3966), .B(n3207), .C(n3967), .D(n3208), .Z(n4146) );
  CANR2X1 U4545 ( .A(n3766), .B(n3203), .C(n5190), .D(n3206), .Z(n4147) );
  CENX1 U4546 ( .A(n4479), .B(n4494), .Z(n3795) );
  CENX1 U4547 ( .A(n4479), .B(n5036), .Z(n3823) );
  CENX1 U4548 ( .A(n4479), .B(n4499), .Z(n3814) );
  CENX1 U4549 ( .A(n4479), .B(n5035), .Z(n3818) );
  CENX1 U4550 ( .A(n4479), .B(n4530), .Z(n3799) );
  CENX1 U4551 ( .A(n4479), .B(n4509), .Z(n3827) );
  CEOX1 U4552 ( .A(n4279), .B(D[31]), .Z(n3763) );
  CEOX1 U4553 ( .A(opera1_copydiv[31]), .B(\intadd_0/n1 ), .Z(n4279) );
  CEOX1 U4554 ( .A(n4274), .B(D[31]), .Z(n3759) );
  CENX1 U4555 ( .A(n3390), .B(\intadd_1/n1 ), .Z(n4274) );
  COND3X1 U4556 ( .A(n4143), .B(n3205), .C(n4264), .D(n4265), .Z(n1495) );
  CND2X1 U4557 ( .A(result_not[59]), .B(n4168), .Z(n4264) );
  CANR2X1 U4558 ( .A(\intadd_1/SUM[26] ), .B(n4484), .C(n4177), .D(n3211), .Z(
        n4265) );
  COND3X1 U4559 ( .A(n4143), .B(n3203), .C(n4268), .D(n4269), .Z(n1493) );
  CND2X1 U4560 ( .A(result_not[61]), .B(n4168), .Z(n4268) );
  CANR2X1 U4561 ( .A(\intadd_1/SUM[28] ), .B(n4484), .C(n4177), .D(n3397), .Z(
        n4269) );
  CENX1 U4562 ( .A(n4478), .B(n4708), .Z(n3780) );
  CNR3XL U4563 ( .A(n5157), .B(n1770), .C(n3201), .Z(n3779) );
  COND3X1 U4564 ( .A(n3465), .B(n5184), .C(n4403), .D(n4404), .Z(n1448) );
  CND2X1 U4565 ( .A(result[42]), .B(n3078), .Z(n4404) );
  COND3X1 U4566 ( .A(result_not[42]), .B(n3323), .C(n4405), .D(n4475), .Z(
        n4403) );
  COND3X1 U4567 ( .A(n3261), .B(n5184), .C(n4394), .D(n4395), .Z(n1451) );
  CND2X1 U4568 ( .A(result[39]), .B(n3078), .Z(n4395) );
  COND3X1 U4569 ( .A(n3326), .B(result_not[39]), .C(n4396), .D(n4475), .Z(
        n4394) );
  CND2X1 U4570 ( .A(result_not[0]), .B(n4168), .Z(n4175) );
  CANR2X1 U4571 ( .A(n4484), .B(n3206), .C(n4177), .D(n335), .Z(n4176) );
  COND3X1 U4572 ( .A(n3453), .B(n5184), .C(n4415), .D(n4416), .Z(n1444) );
  CND2X1 U4573 ( .A(result[46]), .B(n3078), .Z(n4416) );
  COND3X1 U4574 ( .A(result_not[46]), .B(n3319), .C(n4417), .D(n5183), .Z(
        n4415) );
  COND3X1 U4575 ( .A(n3464), .B(n5184), .C(n4409), .D(n4410), .Z(n1446) );
  CND2X1 U4576 ( .A(result[44]), .B(n3078), .Z(n4410) );
  COND3X1 U4577 ( .A(result_not[44]), .B(n3321), .C(n4411), .D(n4475), .Z(
        n4409) );
  COND3X1 U4578 ( .A(n3466), .B(n5184), .C(n4397), .D(n4398), .Z(n1450) );
  CND2X1 U4579 ( .A(result[40]), .B(n3078), .Z(n4398) );
  COND3X1 U4580 ( .A(result_not[40]), .B(n3325), .C(n4399), .D(n5183), .Z(
        n4397) );
  COND3X1 U4581 ( .A(n3478), .B(n5184), .C(n4391), .D(n4392), .Z(n1452) );
  CND2X1 U4582 ( .A(result[38]), .B(n3078), .Z(n4392) );
  COND3X1 U4583 ( .A(result_not[38]), .B(n3327), .C(n4393), .D(n4475), .Z(
        n4391) );
  COND3X1 U4584 ( .A(n3246), .B(n5184), .C(n4412), .D(n4413), .Z(n1445) );
  CND2X1 U4585 ( .A(result[45]), .B(n3078), .Z(n4413) );
  COND3X1 U4586 ( .A(n3320), .B(result_not[45]), .C(n4414), .D(n5183), .Z(
        n4412) );
  COND3X1 U4587 ( .A(n3251), .B(n5184), .C(n4406), .D(n4407), .Z(n1447) );
  CND2X1 U4588 ( .A(result[43]), .B(n3078), .Z(n4407) );
  COND3X1 U4589 ( .A(n3322), .B(result_not[43]), .C(n4408), .D(n4475), .Z(
        n4406) );
  COND3X1 U4590 ( .A(n3256), .B(n4281), .C(n4400), .D(n4401), .Z(n1449) );
  CND2X1 U4591 ( .A(result[41]), .B(n3078), .Z(n4401) );
  COND3X1 U4592 ( .A(n3324), .B(result_not[41]), .C(n4402), .D(n4475), .Z(
        n4400) );
  CND2X1 U4593 ( .A(result_not[63]), .B(n5186), .Z(n4272) );
  CANR2X1 U4594 ( .A(n3958), .B(n3759), .C(n4177), .D(n3396), .Z(n4273) );
  COND3X1 U4595 ( .A(n4143), .B(n3202), .C(n4270), .D(n4271), .Z(n1492) );
  CND2X1 U4596 ( .A(result_not[62]), .B(n5186), .Z(n4270) );
  CANR2X1 U4597 ( .A(\intadd_1/SUM[29] ), .B(n4484), .C(n4177), .D(n3393), .Z(
        n4271) );
  COND3X1 U4598 ( .A(n4143), .B(n3204), .C(n4266), .D(n4267), .Z(n1494) );
  CND2X1 U4599 ( .A(result_not[60]), .B(n5186), .Z(n4266) );
  CANR2X1 U4600 ( .A(\intadd_1/SUM[27] ), .B(n4484), .C(n4177), .D(n3391), .Z(
        n4267) );
  CND2X1 U4601 ( .A(D[0]), .B(opera1_copy[0]), .Z(\intadd_1/CI ) );
  CANR4CX1 U4602 ( .A(n3201), .B(n3758), .C(n4482), .D(n1770), .Z(n3756) );
  CND4X1 U4603 ( .A(n4059), .B(n4060), .C(n4061), .D(n4062), .Z(n1571) );
  CANR2X1 U4604 ( .A(n5188), .B(D[18]), .C(n1803), .D(n5191), .Z(n4060) );
  CANR2X1 U4605 ( .A(n5187), .B(n3233), .C(n3958), .D(n3235), .Z(n4059) );
  CANR2X1 U4606 ( .A(n5178), .B(n3237), .C(n5190), .D(n3234), .Z(n4061) );
  CND4X1 U4607 ( .A(n4072), .B(n4073), .C(n4074), .D(n4075), .Z(n1569) );
  CANR2X1 U4608 ( .A(n5188), .B(D[20]), .C(n1804), .D(n3753), .Z(n4073) );
  CANR2X1 U4609 ( .A(n5187), .B(n3228), .C(n3958), .D(n3230), .Z(n4072) );
  CANR2X1 U4610 ( .A(n5178), .B(n3232), .C(n5190), .D(n3229), .Z(n4074) );
  CND4X1 U4611 ( .A(n4085), .B(n4086), .C(n4087), .D(n4088), .Z(n1567) );
  CANR2X1 U4612 ( .A(n5188), .B(D[22]), .C(n1805), .D(n5191), .Z(n4086) );
  CANR2X1 U4613 ( .A(n5187), .B(n3223), .C(n5177), .D(n3225), .Z(n4085) );
  CANR2X1 U4614 ( .A(n5178), .B(n3227), .C(n5190), .D(n3224), .Z(n4087) );
  CND4X1 U4615 ( .A(n4098), .B(n4099), .C(n4100), .D(n4101), .Z(n1565) );
  CANR2X1 U4616 ( .A(n5188), .B(D[24]), .C(n1806), .D(n3753), .Z(n4099) );
  CANR2X1 U4617 ( .A(n5187), .B(n3218), .C(n3958), .D(n3220), .Z(n4098) );
  CANR2X1 U4618 ( .A(n5178), .B(n3222), .C(n5190), .D(n3219), .Z(n4100) );
  CND4X1 U4619 ( .A(n4111), .B(n4112), .C(n4113), .D(n4114), .Z(n1563) );
  CANR2X1 U4620 ( .A(n5188), .B(D[26]), .C(n1807), .D(n5191), .Z(n4112) );
  CANR2X1 U4621 ( .A(n5187), .B(n3213), .C(n4484), .D(n3215), .Z(n4111) );
  CANR2X1 U4622 ( .A(n5178), .B(n3217), .C(n5190), .D(n3214), .Z(n4113) );
  CND4X1 U4623 ( .A(n4124), .B(n4125), .C(n4126), .D(n4127), .Z(n1561) );
  CANR2X1 U4624 ( .A(n5188), .B(D[28]), .C(n1808), .D(n5191), .Z(n4125) );
  CANR2X1 U4625 ( .A(n5187), .B(n3205), .C(n5177), .D(n3210), .Z(n4124) );
  CANR2X1 U4626 ( .A(n5178), .B(n3212), .C(n5190), .D(n3209), .Z(n4126) );
  CND4X1 U4627 ( .A(n4065), .B(n4066), .C(n4067), .D(n4853), .Z(n1570) );
  CANR2X1 U4628 ( .A(n3967), .B(n3235), .C(n1804), .D(n5188), .Z(n4066) );
  CANR2X1 U4629 ( .A(n3949), .B(n3232), .C(n4483), .D(D[18]), .Z(n4065) );
  CANR2X1 U4630 ( .A(n5190), .B(n3230), .C(n3966), .D(n3234), .Z(n4067) );
  CND4X1 U4631 ( .A(n4091), .B(n4092), .C(n4093), .D(n4806), .Z(n1566) );
  CANR2X1 U4632 ( .A(n3967), .B(n3225), .C(n1806), .D(n5188), .Z(n4092) );
  CANR2X1 U4633 ( .A(n3949), .B(n3222), .C(n4483), .D(D[22]), .Z(n4091) );
  CANR2X1 U4634 ( .A(n5190), .B(n3220), .C(n3966), .D(n3224), .Z(n4093) );
  CND4X1 U4635 ( .A(n4117), .B(n4118), .C(n4119), .D(n4802), .Z(n1562) );
  CANR2X1 U4636 ( .A(n3967), .B(n3215), .C(n1808), .D(n5188), .Z(n4118) );
  CANR2X1 U4637 ( .A(n3949), .B(n3212), .C(n4483), .D(D[26]), .Z(n4117) );
  CANR2X1 U4638 ( .A(n5190), .B(n3210), .C(n3966), .D(n3214), .Z(n4119) );
  CANR3X1 U4639 ( .A(n4483), .B(n4488), .C(n3166), .D(n3771), .Z(n3770) );
  CANR11X1 U4640 ( .A(n3179), .B(cin2a), .C(n5181), .D(n3779), .Z(n3768) );
  CND2X1 U4641 ( .A(D[0]), .B(opera1_copydiv[0]), .Z(\intadd_0/CI ) );
  CNR2IX1 U4642 ( .B(cin1a), .A(n3644), .Z(n3635) );
  CEOX1 U4643 ( .A(n3136), .B(n4984), .Z(n3644) );
  COND3X1 U4644 ( .A(n4952), .B(n3162), .C(n3126), .D(n3626), .Z(n3616) );
  CANR2X1 U4645 ( .A(n3136), .B(n3162), .C(n4952), .D(n4986), .Z(n3626) );
  COND3X1 U4646 ( .A(n4920), .B(n3159), .C(n3101), .D(n3606), .Z(n3596) );
  CANR2X1 U4647 ( .A(n3136), .B(n3159), .C(n4920), .D(n4986), .Z(n3606) );
  COND3X1 U4648 ( .A(n3136), .B(n3155), .C(n3098), .D(n3586), .Z(n3576) );
  CANR2X1 U4649 ( .A(n3156), .B(n3136), .C(n4928), .D(n3155), .Z(n3586) );
  COND3X1 U4650 ( .A(n3136), .B(n3151), .C(n3096), .D(n3566), .Z(n3556) );
  CANR2X1 U4651 ( .A(n3152), .B(n3136), .C(n4876), .D(n3151), .Z(n3566) );
  COND3X1 U4652 ( .A(n3136), .B(n3147), .C(n3094), .D(n3546), .Z(n3533) );
  CANR2X1 U4653 ( .A(n3148), .B(n3136), .C(n4870), .D(n3147), .Z(n3546) );
  COND3X1 U4654 ( .A(n3136), .B(n3143), .C(n3092), .D(n3525), .Z(n3513) );
  CANR2X1 U4655 ( .A(n3144), .B(n3136), .C(n4818), .D(n3143), .Z(n3525) );
  COND3X1 U4656 ( .A(n3136), .B(n3141), .C(n3091), .D(n3515), .Z(n3501) );
  CANR2X1 U4657 ( .A(n3142), .B(n3136), .C(n4812), .D(n3141), .Z(n3515) );
  COND3X1 U4658 ( .A(n3136), .B(n3145), .C(n3093), .D(n3535), .Z(n3523) );
  CANR2X1 U4659 ( .A(n3146), .B(n3136), .C(n4817), .D(n3145), .Z(n3535) );
  CNR2X1 U4660 ( .A(n3497), .B(n4694), .Z(n3487) );
  COND3X1 U4661 ( .A(n3136), .B(n3163), .C(n3635), .D(n3636), .Z(n3625) );
  CANR2X1 U4662 ( .A(n3164), .B(n3136), .C(n4972), .D(n3163), .Z(n3636) );
  COND3X1 U4663 ( .A(n3136), .B(n3160), .C(n3102), .D(n3615), .Z(n3605) );
  CANR2X1 U4664 ( .A(n3136), .B(n4967), .C(n4969), .D(n3160), .Z(n3615) );
  COND3X1 U4665 ( .A(n3136), .B(n3157), .C(n3099), .D(n3595), .Z(n3585) );
  CANR2X1 U4666 ( .A(n4921), .B(n3157), .C(n3136), .D(n3158), .Z(n3595) );
  COND3X1 U4667 ( .A(n3136), .B(n3153), .C(n3097), .D(n3575), .Z(n3565) );
  CANR2X1 U4668 ( .A(n4862), .B(n3136), .C(n4863), .D(n3153), .Z(n3575) );
  COND3X1 U4669 ( .A(n3136), .B(n3149), .C(n3095), .D(n3555), .Z(n3544) );
  CANR2X1 U4670 ( .A(n4866), .B(n3136), .C(n4868), .D(n3149), .Z(n3555) );
  CND2X1 U4671 ( .A(n3504), .B(n3090), .Z(n3497) );
  CANR4CX1 U4672 ( .A(n4986), .B(n3140), .C(n4571), .D(n3505), .Z(n3504) );
  CANR1XL U4673 ( .A(n4986), .B(n3140), .C(n4697), .Z(n3505) );
  CNR2X1 U4674 ( .A(n4478), .B(n5074), .Z(n3891) );
  CNR2X1 U4675 ( .A(n4478), .B(n5052), .Z(n3849) );
  CNR2X1 U4676 ( .A(n4478), .B(n5063), .Z(n3870) );
  COND3X1 U4677 ( .A(n4143), .B(n3223), .C(n4252), .D(n4253), .Z(n1501) );
  CND2X1 U4678 ( .A(result_not[53]), .B(n4168), .Z(n4252) );
  CANR2X1 U4679 ( .A(\intadd_1/SUM[20] ), .B(n4484), .C(n4177), .D(n3226), .Z(
        n4253) );
  COND3X1 U4680 ( .A(n4143), .B(n3218), .C(n4256), .D(n4257), .Z(n1499) );
  CND2X1 U4681 ( .A(result_not[55]), .B(n4168), .Z(n4256) );
  CANR2X1 U4682 ( .A(\intadd_1/SUM[22] ), .B(n4484), .C(n4177), .D(n3221), .Z(
        n4257) );
  COND3X1 U4683 ( .A(n4143), .B(n3213), .C(n4260), .D(n4261), .Z(n1497) );
  CND2X1 U4684 ( .A(result_not[57]), .B(n4168), .Z(n4260) );
  CANR2X1 U4685 ( .A(\intadd_1/SUM[24] ), .B(n4484), .C(n4177), .D(n3216), .Z(
        n4261) );
  CND3XL U4686 ( .A(n5192), .B(n3137), .C(n3487), .Z(n3485) );
  CND3XL U4687 ( .A(n3488), .B(n3489), .C(n4690), .Z(n3484) );
  COND3X1 U4688 ( .A(n4143), .B(n3212), .C(n4262), .D(n4263), .Z(n1496) );
  CND2X1 U4689 ( .A(result_not[58]), .B(n5186), .Z(n4262) );
  CANR2X1 U4690 ( .A(\intadd_1/SUM[25] ), .B(n4484), .C(n4177), .D(n3392), .Z(
        n4263) );
  COND3X1 U4691 ( .A(n4143), .B(n3217), .C(n4258), .D(n4259), .Z(n1498) );
  CND2X1 U4692 ( .A(result_not[56]), .B(n5186), .Z(n4258) );
  CANR2X1 U4693 ( .A(\intadd_1/SUM[23] ), .B(n4484), .C(n4177), .D(n3423), .Z(
        n4259) );
  COND3X1 U4694 ( .A(n4143), .B(n3222), .C(n4254), .D(n4255), .Z(n1500) );
  CND2X1 U4695 ( .A(result_not[54]), .B(n5186), .Z(n4254) );
  CANR2X1 U4696 ( .A(\intadd_1/SUM[21] ), .B(n4484), .C(n4177), .D(n3424), .Z(
        n4255) );
  COND4CX1 U4697 ( .A(n3497), .B(n3138), .C(n3489), .D(n5192), .Z(n3495) );
  CANR2X1 U4698 ( .A(n4694), .B(n3494), .C(n4476), .D(opera1_copy[29]), .Z(
        n3496) );
  CND3XL U4699 ( .A(n3497), .B(n3139), .C(n3500), .Z(n3499) );
  COND4CX1 U4700 ( .A(n3502), .B(n4477), .C(n3494), .D(n4571), .Z(n3498) );
  COND11X1 U4701 ( .A(n3127), .B(n3140), .C(n3501), .D(n4486), .Z(n3500) );
  CNR2X1 U4702 ( .A(n3084), .B(n4486), .Z(n3493) );
  COND3X1 U4703 ( .A(n1741), .B(n5184), .C(n4385), .D(n4386), .Z(n1454) );
  CND2X1 U4704 ( .A(result[36]), .B(n3078), .Z(n4386) );
  COND3X1 U4705 ( .A(result_not[36]), .B(n3329), .C(n4387), .D(n4309), .Z(
        n4385) );
  COND3X1 U4706 ( .A(n3477), .B(n5184), .C(n4379), .D(n4380), .Z(n1456) );
  CND2X1 U4707 ( .A(result[34]), .B(n3078), .Z(n4380) );
  COND3X1 U4708 ( .A(result_not[34]), .B(n3331), .C(n4381), .D(n5183), .Z(
        n4379) );
  COND3X1 U4709 ( .A(n3482), .B(n5184), .C(n4373), .D(n4374), .Z(n1458) );
  CND2X1 U4710 ( .A(result[32]), .B(n3078), .Z(n4374) );
  COND3X1 U4711 ( .A(result_not[32]), .B(n3333), .C(n4375), .D(n5183), .Z(
        n4373) );
  COND3X1 U4712 ( .A(n3373), .B(n5184), .C(n4367), .D(n4368), .Z(n1460) );
  CND2X1 U4713 ( .A(result[30]), .B(n3078), .Z(n4368) );
  COND3X1 U4714 ( .A(result_not[30]), .B(n3335), .C(n4369), .D(n4475), .Z(
        n4367) );
  COND3X1 U4715 ( .A(n3266), .B(n5184), .C(n4388), .D(n4389), .Z(n1453) );
  CND2X1 U4716 ( .A(result[37]), .B(n3078), .Z(n4389) );
  COND3X1 U4717 ( .A(n3328), .B(result_not[37]), .C(n4390), .D(n4475), .Z(
        n4388) );
  COND3X1 U4718 ( .A(n3272), .B(n5184), .C(n4382), .D(n4383), .Z(n1455) );
  CND2X1 U4719 ( .A(result[35]), .B(n3078), .Z(n4383) );
  COND3X1 U4720 ( .A(n3330), .B(result_not[35]), .C(n4384), .D(n4309), .Z(
        n4382) );
  COND3X1 U4721 ( .A(n3316), .B(n5184), .C(n4376), .D(n4377), .Z(n1457) );
  CND2X1 U4722 ( .A(result[33]), .B(n3078), .Z(n4377) );
  COND3X1 U4723 ( .A(n3332), .B(result_not[33]), .C(n4378), .D(n4309), .Z(
        n4376) );
  COND3X1 U4724 ( .A(n3284), .B(n5184), .C(n4370), .D(n4371), .Z(n1459) );
  CND2X1 U4725 ( .A(result[31]), .B(n3078), .Z(n4371) );
  COND3X1 U4726 ( .A(n3334), .B(result_not[31]), .C(n4372), .D(n5183), .Z(
        n4370) );
  COND2X1 U4727 ( .A(\intadd_1/SUM[3] ), .B(n3276), .C(\intadd_1/SUM[4] ), .D(
        n4487), .Z(n3977) );
  COND2X1 U4728 ( .A(n4485), .B(n3266), .C(\intadd_1/SUM[2] ), .D(n3277), .Z(
        n3974) );
  COND2X1 U4729 ( .A(n1741), .B(n4482), .C(\intadd_0/SUM[3] ), .D(n3275), .Z(
        n3975) );
  CND4X1 U4730 ( .A(n3981), .B(n3982), .C(n3983), .D(n3984), .Z(n1583) );
  CANR2X1 U4731 ( .A(n5187), .B(n3263), .C(n4484), .D(n3265), .Z(n3981) );
  CANR2X1 U4732 ( .A(n5188), .B(D[6]), .C(n1797), .D(n4483), .Z(n3982) );
  CANR2X1 U4733 ( .A(n5178), .B(n3267), .C(n5190), .D(n3264), .Z(n3983) );
  CND4X1 U4734 ( .A(n3994), .B(n3995), .C(n3996), .D(n3997), .Z(n1581) );
  CANR2X1 U4735 ( .A(n5187), .B(n3258), .C(n5177), .D(n3260), .Z(n3994) );
  CANR2X1 U4736 ( .A(n5188), .B(D[8]), .C(n1798), .D(n4483), .Z(n3995) );
  CANR2X1 U4737 ( .A(n5178), .B(n3262), .C(n5190), .D(n3259), .Z(n3996) );
  CND4X1 U4738 ( .A(n4007), .B(n4008), .C(n4009), .D(n4010), .Z(n1579) );
  CANR2X1 U4739 ( .A(n5187), .B(n3253), .C(n5177), .D(n3255), .Z(n4007) );
  CANR2X1 U4740 ( .A(n5188), .B(D[10]), .C(n1799), .D(n5191), .Z(n4008) );
  CANR2X1 U4741 ( .A(n5178), .B(n3257), .C(n5190), .D(n3254), .Z(n4009) );
  CND4X1 U4742 ( .A(n4020), .B(n4021), .C(n4022), .D(n4023), .Z(n1577) );
  CANR2X1 U4743 ( .A(n5187), .B(n3248), .C(n3958), .D(n3250), .Z(n4020) );
  CANR2X1 U4744 ( .A(n5188), .B(D[12]), .C(n1800), .D(n5191), .Z(n4021) );
  CANR2X1 U4745 ( .A(n5178), .B(n3252), .C(n5190), .D(n3249), .Z(n4022) );
  CND4X1 U4746 ( .A(n4033), .B(n4034), .C(n4035), .D(n4036), .Z(n1575) );
  CANR2X1 U4747 ( .A(n5188), .B(D[14]), .C(n1801), .D(n4483), .Z(n4034) );
  CANR2X1 U4748 ( .A(n5187), .B(n3243), .C(n3958), .D(n3245), .Z(n4033) );
  CANR2X1 U4749 ( .A(n5178), .B(n3247), .C(n5190), .D(n3244), .Z(n4035) );
  CND4X1 U4750 ( .A(n4046), .B(n4047), .C(n4048), .D(n4049), .Z(n1573) );
  CANR2X1 U4751 ( .A(n5188), .B(D[16]), .C(n1802), .D(n5191), .Z(n4047) );
  CANR2X1 U4752 ( .A(n5187), .B(n3238), .C(n3958), .D(n3240), .Z(n4046) );
  CANR2X1 U4753 ( .A(n5178), .B(n3242), .C(n5190), .D(n3239), .Z(n4048) );
  CND4X1 U4754 ( .A(n3987), .B(n3988), .C(n3989), .D(n4962), .Z(n1582) );
  CANR2X1 U4755 ( .A(n3949), .B(n3262), .C(n5191), .D(D[6]), .Z(n3987) );
  CANR2X1 U4756 ( .A(n5190), .B(n3260), .C(n3966), .D(n3264), .Z(n3989) );
  CANR2X1 U4757 ( .A(n3967), .B(n3265), .C(n1798), .D(n5188), .Z(n3988) );
  CND4X1 U4758 ( .A(n4013), .B(n4014), .C(n4015), .D(n4914), .Z(n1578) );
  CANR2X1 U4759 ( .A(n3949), .B(n3252), .C(n5191), .D(D[10]), .Z(n4013) );
  CANR2X1 U4760 ( .A(n5190), .B(n3250), .C(n3966), .D(n3254), .Z(n4015) );
  CANR2X1 U4761 ( .A(n3967), .B(n3255), .C(n1800), .D(n5188), .Z(n4014) );
  CND4X1 U4762 ( .A(n4039), .B(n4040), .C(n4041), .D(n4857), .Z(n1574) );
  CANR2X1 U4763 ( .A(n3967), .B(n3245), .C(n1802), .D(n5188), .Z(n4040) );
  CANR2X1 U4764 ( .A(n3949), .B(n3242), .C(n5191), .D(D[14]), .Z(n4039) );
  CANR2X1 U4765 ( .A(n5190), .B(n3240), .C(n3966), .D(n3244), .Z(n4041) );
  CENX1 U4766 ( .A(n4479), .B(n5101), .Z(n3937) );
  CANR1XL U4767 ( .A(n3091), .B(muordi), .C(n3104), .Z(n3519) );
  CENX1 U4768 ( .A(n4986), .B(n4952), .Z(n3659) );
  COND3X1 U4769 ( .A(n4143), .B(n3238), .C(n4240), .D(n4241), .Z(n1507) );
  CND2X1 U4770 ( .A(result_not[47]), .B(n4168), .Z(n4240) );
  CANR2X1 U4771 ( .A(\intadd_1/SUM[14] ), .B(n5177), .C(n4177), .D(n3241), .Z(
        n4241) );
  CANR11X1 U4772 ( .A(n3094), .B(n4870), .C(n3492), .D(n5192), .Z(n3543) );
  CENX1 U4773 ( .A(n3136), .B(n4923), .Z(n3668) );
  CENX1 U4774 ( .A(n3136), .B(n4971), .Z(n3652) );
  COND3X1 U4775 ( .A(n4482), .B(n3284), .C(n3933), .D(n3934), .Z(n1589) );
  CANR2X1 U4776 ( .A(n5188), .B(D[0]), .C(result_copy[30]), .D(n5189), .Z(
        n3933) );
  CANR1XL U4777 ( .A(n5190), .B(n3476), .C(n3935), .Z(n3934) );
  CANR11X1 U4778 ( .A(n3169), .B(n3916), .C(n3778), .D(n3922), .Z(n3921) );
  CAN2X1 U4779 ( .A(n4519), .B(n3775), .Z(n3922) );
  CANR11X1 U4780 ( .A(n3168), .B(n3926), .C(n3778), .D(n3932), .Z(n3931) );
  CAN2X1 U4781 ( .A(n4528), .B(n3775), .Z(n3932) );
  CANR11X1 U4782 ( .A(n3170), .B(n3905), .C(n5181), .D(n3911), .Z(n3910) );
  CAN2X1 U4783 ( .A(n4501), .B(n3775), .Z(n3911) );
  CNR2X1 U4784 ( .A(n4478), .B(n5085), .Z(n3912) );
  CNR2X1 U4785 ( .A(n4818), .B(n3523), .Z(n3524) );
  CNR2X1 U4786 ( .A(n4817), .B(n3533), .Z(n3534) );
  CNR2X1 U4787 ( .A(n4812), .B(n3513), .Z(n3514) );
  CNR2X1 U4788 ( .A(n4700), .B(n3501), .Z(n3502) );
  COND2X1 U4789 ( .A(n4481), .B(\intadd_0/B[22] ), .C(n4480), .D(n3711), .Z(
        n1663) );
  CENX1 U4790 ( .A(n3710), .B(n3712), .Z(n3711) );
  CND2X1 U4791 ( .A(cin1b), .B(n3644), .Z(n3650) );
  COND1XL U4792 ( .A(n4481), .B(\intadd_0/B[24] ), .C(n3716), .Z(n1661) );
  COND3X1 U4793 ( .A(n3110), .B(n3717), .C(n3718), .D(n4481), .Z(n3716) );
  COND3X1 U4794 ( .A(n4143), .B(n3233), .C(n4244), .D(n4245), .Z(n1505) );
  CND2X1 U4795 ( .A(result_not[49]), .B(n4168), .Z(n4244) );
  CANR2X1 U4796 ( .A(\intadd_1/SUM[16] ), .B(n3958), .C(n4177), .D(n3236), .Z(
        n4245) );
  COND3X1 U4797 ( .A(n4143), .B(n3228), .C(n4248), .D(n4249), .Z(n1503) );
  CND2X1 U4798 ( .A(result_not[51]), .B(n4168), .Z(n4248) );
  CANR2X1 U4799 ( .A(\intadd_1/SUM[18] ), .B(n4484), .C(n4177), .D(n3231), .Z(
        n4249) );
  COND3X1 U4800 ( .A(n3772), .B(n3373), .C(n3923), .D(n3924), .Z(n1591) );
  CANR2X1 U4801 ( .A(result_copy[28]), .B(n5189), .C(result_copy[29]), .D(
        n4483), .Z(n3924) );
  CENX1 U4802 ( .A(n3926), .B(n3920), .Z(n3925) );
  COND3X1 U4803 ( .A(n3772), .B(n3366), .C(n3902), .D(n3903), .Z(n1595) );
  CANR2X1 U4804 ( .A(result_copy[24]), .B(n5189), .C(result_copy[25]), .D(
        n4483), .Z(n3903) );
  CENX1 U4805 ( .A(n3905), .B(n3899), .Z(n3904) );
  COND3X1 U4806 ( .A(n3772), .B(n3376), .C(n3913), .D(n3914), .Z(n1593) );
  CANR2X1 U4807 ( .A(result_copy[26]), .B(n5189), .C(result_copy[27]), .D(
        n4483), .Z(n3914) );
  CENX1 U4808 ( .A(n3909), .B(n3916), .Z(n3915) );
  COND3X1 U4809 ( .A(n4482), .B(n3482), .C(n3939), .D(n4990), .Z(n1588) );
  CANR2X1 U4810 ( .A(n1773), .B(n5188), .C(n3948), .D(n3949), .Z(n3939) );
  CANR3X1 U4811 ( .A(n4991), .B(n4481), .C(n3942), .D(n3943), .Z(n3940) );
  CNR3XL U4812 ( .A(n3284), .B(n3944), .C(n5157), .Z(n3943) );
  COND4CX1 U4813 ( .A(n5192), .B(n3544), .C(n3549), .D(n3148), .Z(n3548) );
  COND4CX1 U4814 ( .A(n5192), .B(n3094), .C(n3550), .D(n4870), .Z(n3547) );
  CNR2X1 U4815 ( .A(n3544), .B(n3103), .Z(n3549) );
  COND4CX1 U4816 ( .A(n5192), .B(n3523), .C(n3528), .D(n3144), .Z(n3527) );
  COND4CX1 U4817 ( .A(n5192), .B(n3092), .C(n3529), .D(n4818), .Z(n3526) );
  CNR2X1 U4818 ( .A(n3523), .B(n3103), .Z(n3528) );
  CND3XL U4819 ( .A(n3513), .B(n3143), .C(n3522), .Z(n3521) );
  COND4CX1 U4820 ( .A(n3524), .B(n4477), .C(n3519), .D(n4728), .Z(n3520) );
  COND11X1 U4821 ( .A(n3127), .B(n3144), .C(n3523), .D(n4486), .Z(n3522) );
  CND3XL U4822 ( .A(n3523), .B(n3145), .C(n3532), .Z(n3531) );
  COND4CX1 U4823 ( .A(n3534), .B(n4477), .C(n3529), .D(n4720), .Z(n3530) );
  COND11X1 U4824 ( .A(n3127), .B(n4815), .C(n3533), .D(n4486), .Z(n3532) );
  COND3X1 U4825 ( .A(n4143), .B(n3227), .C(n4250), .D(n4251), .Z(n1502) );
  CND2X1 U4826 ( .A(result_not[52]), .B(n4168), .Z(n4250) );
  CANR2X1 U4827 ( .A(\intadd_1/SUM[19] ), .B(n4484), .C(n4177), .D(n3426), .Z(
        n4251) );
  COND3X1 U4828 ( .A(n4143), .B(n3232), .C(n4246), .D(n4247), .Z(n1504) );
  CND2X1 U4829 ( .A(result_not[50]), .B(n4168), .Z(n4246) );
  CANR2X1 U4830 ( .A(\intadd_1/SUM[17] ), .B(n4484), .C(n4177), .D(n3451), .Z(
        n4247) );
  COND3X1 U4831 ( .A(n4143), .B(n3237), .C(n4242), .D(n4243), .Z(n1506) );
  CND2X1 U4832 ( .A(result_not[48]), .B(n4168), .Z(n4242) );
  CANR2X1 U4833 ( .A(\intadd_1/SUM[15] ), .B(n5177), .C(n4177), .D(n3452), .Z(
        n4243) );
  COND3X1 U4834 ( .A(n4143), .B(n3242), .C(n4238), .D(n4239), .Z(n1508) );
  CND2X1 U4835 ( .A(result_not[46]), .B(n4168), .Z(n4238) );
  CANR2X1 U4836 ( .A(\intadd_1/SUM[13] ), .B(n4484), .C(n4177), .D(n3453), .Z(
        n4239) );
  COND4CX1 U4837 ( .A(n5192), .B(n3501), .C(n3508), .D(n3140), .Z(n3507) );
  COND4CX1 U4838 ( .A(n5192), .B(n3090), .C(n3509), .D(n4700), .Z(n3506) );
  CNR2X1 U4839 ( .A(n3501), .B(n3103), .Z(n3508) );
  COND4CX1 U4840 ( .A(n5192), .B(n3513), .C(n3518), .D(n3142), .Z(n3517) );
  COND4CX1 U4841 ( .A(n5192), .B(n3091), .C(n3519), .D(n4812), .Z(n3516) );
  CNR2X1 U4842 ( .A(n3513), .B(n3103), .Z(n3518) );
  COND3X1 U4843 ( .A(n3512), .B(n5192), .C(n3501), .D(n3141), .Z(n3511) );
  COND4CX1 U4844 ( .A(n3514), .B(n4477), .C(n3509), .D(n4568), .Z(n3510) );
  CNR3XL U4845 ( .A(n3127), .B(n3142), .C(n3513), .Z(n3512) );
  COND3X1 U4846 ( .A(n3375), .B(n4281), .C(n4343), .D(n4344), .Z(n1468) );
  CND2X1 U4847 ( .A(result[22]), .B(n3078), .Z(n4344) );
  COND3X1 U4848 ( .A(result_not[22]), .B(n3343), .C(n4345), .D(n5183), .Z(
        n4343) );
  COND3X1 U4849 ( .A(n3369), .B(n4281), .C(n4349), .D(n4350), .Z(n1466) );
  CND2X1 U4850 ( .A(result[24]), .B(n3078), .Z(n4350) );
  COND3X1 U4851 ( .A(result_not[24]), .B(n3341), .C(n4351), .D(n4475), .Z(
        n4349) );
  COND3X1 U4852 ( .A(n3366), .B(n5184), .C(n4355), .D(n4356), .Z(n1464) );
  CND2X1 U4853 ( .A(result[26]), .B(n3078), .Z(n4356) );
  COND3X1 U4854 ( .A(result_not[26]), .B(n3339), .C(n4357), .D(n5183), .Z(
        n4355) );
  COND3X1 U4855 ( .A(n3376), .B(n5184), .C(n4361), .D(n4362), .Z(n1462) );
  CND2X1 U4856 ( .A(result[28]), .B(n3078), .Z(n4362) );
  COND3X1 U4857 ( .A(result_not[28]), .B(n3337), .C(n4363), .D(n4475), .Z(
        n4361) );
  COND3X1 U4858 ( .A(n3294), .B(n5184), .C(n4340), .D(n4341), .Z(n1469) );
  CND2X1 U4859 ( .A(result[21]), .B(n3078), .Z(n4341) );
  COND3X1 U4860 ( .A(n3344), .B(result_not[21]), .C(n4342), .D(n4309), .Z(
        n4340) );
  COND3X1 U4861 ( .A(n3296), .B(n5184), .C(n4346), .D(n4347), .Z(n1467) );
  CND2X1 U4862 ( .A(result[23]), .B(n3078), .Z(n4347) );
  COND3X1 U4863 ( .A(n3342), .B(result_not[23]), .C(n4348), .D(n4475), .Z(
        n4346) );
  COND3X1 U4864 ( .A(n3286), .B(n5184), .C(n4352), .D(n4353), .Z(n1465) );
  CND2X1 U4865 ( .A(result[25]), .B(n3078), .Z(n4353) );
  COND3X1 U4866 ( .A(n3340), .B(result_not[25]), .C(n4354), .D(n4475), .Z(
        n4352) );
  COND3X1 U4867 ( .A(n3285), .B(n5184), .C(n4358), .D(n4359), .Z(n1463) );
  CND2X1 U4868 ( .A(result[27]), .B(n3078), .Z(n4359) );
  COND3X1 U4869 ( .A(n3338), .B(result_not[27]), .C(n4360), .D(n4309), .Z(
        n4358) );
  COND3X1 U4870 ( .A(n3293), .B(n5184), .C(n4364), .D(n4365), .Z(n1461) );
  CND2X1 U4871 ( .A(result[29]), .B(n3078), .Z(n4365) );
  COND3X1 U4872 ( .A(n3336), .B(result_not[29]), .C(n4366), .D(n5183), .Z(
        n4364) );
  CANR2X1 U4873 ( .A(result_copy[27]), .B(n5189), .C(result_copy[28]), .D(
        n4483), .Z(n3918) );
  COND1XL U4874 ( .A(n4519), .B(n3178), .C(n3921), .Z(n3919) );
  COND3X1 U4875 ( .A(n3772), .B(n3284), .C(n3927), .D(n3928), .Z(n1590) );
  CANR2X1 U4876 ( .A(result_copy[29]), .B(n5189), .C(result_copy[30]), .D(
        n4483), .Z(n3928) );
  COND1XL U4877 ( .A(n4528), .B(n3178), .C(n3931), .Z(n3929) );
  COND3X1 U4878 ( .A(n3772), .B(n3285), .C(n3906), .D(n3907), .Z(n1594) );
  CANR2X1 U4879 ( .A(result_copy[25]), .B(n5189), .C(result_copy[26]), .D(
        n4483), .Z(n3907) );
  COND1XL U4880 ( .A(n4501), .B(n3178), .C(n3910), .Z(n3908) );
  COND1XL U4881 ( .A(n4481), .B(\intadd_0/B[26] ), .C(n3722), .Z(n1659) );
  COND3X1 U4882 ( .A(n3108), .B(n3723), .C(n3724), .D(n4481), .Z(n3722) );
  COND1XL U4883 ( .A(n4481), .B(n1772), .C(n3728), .Z(n1657) );
  COND3X1 U4884 ( .A(n3106), .B(n3729), .C(n3730), .D(n4481), .Z(n3728) );
  COND1XL U4885 ( .A(n3441), .B(n4477), .C(n3551), .Z(n243) );
  CANR4CX1 U4886 ( .A(n3552), .B(n3550), .C(n4841), .D(n3553), .Z(n3551) );
  CNR3XL U4887 ( .A(n4476), .B(n4868), .C(n3556), .Z(n3552) );
  CNR3XL U4888 ( .A(n3554), .B(n4841), .C(n3094), .Z(n3553) );
  COND1XL U4889 ( .A(n3405), .B(n4477), .C(n3540), .Z(n245) );
  CANR1XL U4890 ( .A(n4734), .B(n3541), .C(n3542), .Z(n3540) );
  CNR3XL U4891 ( .A(n3543), .B(n4736), .C(n3093), .Z(n3542) );
  COND11X1 U4892 ( .A(n4476), .B(n4870), .C(n3544), .D(n3539), .Z(n3541) );
  CND4X1 U4893 ( .A(n3950), .B(n3951), .C(n3952), .D(n5110), .Z(n1587) );
  CANR2X1 U4894 ( .A(n5187), .B(n3313), .C(n4484), .D(n3315), .Z(n3950) );
  CANR2X1 U4895 ( .A(n5188), .B(D[2]), .C(n1773), .D(n5191), .Z(n3951) );
  CANR2X1 U4896 ( .A(n5178), .B(n3948), .C(n5190), .D(n3314), .Z(n3952) );
  CND4X1 U4897 ( .A(n3959), .B(n3960), .C(n3961), .D(n4958), .Z(n1586) );
  CANR2X1 U4898 ( .A(n3949), .B(n3312), .C(n5191), .D(D[2]), .Z(n3959) );
  CANR2X1 U4899 ( .A(n5190), .B(n3270), .C(n3966), .D(n3314), .Z(n3961) );
  CANR2X1 U4900 ( .A(n3967), .B(n3315), .C(n1796), .D(n5188), .Z(n3960) );
  CANR4CX1 U4901 ( .A(n3730), .B(n3732), .C(n4481), .D(n3734), .Z(n3733) );
  CNR3X1 U4902 ( .A(n3944), .B(n1770), .C(n5157), .Z(n3766) );
  CANR3X1 U4903 ( .A(n4148), .B(n3944), .C(n260), .D(n3479), .Z(n4166) );
  CND4X1 U4904 ( .A(n4174), .B(n3361), .C(i[5]), .D(n4275), .Z(n4148) );
  CENX1 U4905 ( .A(opera2[43]), .B(n4478), .Z(n4025) );
  CENX1 U4906 ( .A(n4986), .B(n4920), .Z(n3670) );
  COND3X1 U4907 ( .A(n3772), .B(n3364), .C(n3787), .D(n3788), .Z(n1618) );
  CANR2X1 U4908 ( .A(result_copy[1]), .B(n5189), .C(result_copy[2]), .D(n5191), 
        .Z(n3788) );
  CANR2X1 U4909 ( .A(result_copy[5]), .B(n5189), .C(result_copy[6]), .D(n3753), 
        .Z(n3806) );
  COND3X1 U4910 ( .A(n3195), .B(n3165), .C(n3809), .D(n3810), .Z(n3807) );
  COND3X1 U4911 ( .A(n4143), .B(n3262), .C(n4222), .D(n4223), .Z(n1516) );
  CND2X1 U4912 ( .A(result_not[38]), .B(n4168), .Z(n4222) );
  CANR2X1 U4913 ( .A(\intadd_1/SUM[5] ), .B(n3958), .C(n4177), .D(n3478), .Z(
        n4223) );
  COND3X1 U4914 ( .A(n4143), .B(n3312), .C(n4214), .D(n4215), .Z(n1520) );
  CND2X1 U4915 ( .A(result_not[34]), .B(n4168), .Z(n4214) );
  CANR2X1 U4916 ( .A(\intadd_1/SUM[1] ), .B(n5177), .C(n4177), .D(n3477), .Z(
        n4215) );
  CND2X1 U4917 ( .A(n3945), .B(n4484), .Z(n4210) );
  CANR2X1 U4918 ( .A(result_not[32]), .B(n4168), .C(n4177), .D(n3482), .Z(
        n4211) );
  CANR2X1 U4919 ( .A(result_copy[10]), .B(n5189), .C(n5191), .D(n3377), .Z(
        n3830) );
  CEOX1 U4920 ( .A(n3828), .B(n3832), .Z(n3831) );
  COND3X1 U4921 ( .A(n3772), .B(n3297), .C(n3843), .D(n3844), .Z(n1606) );
  CANR2X1 U4922 ( .A(result_copy[13]), .B(n5189), .C(result_copy[14]), .D(
        n4483), .Z(n3844) );
  COND3X1 U4923 ( .A(n3192), .B(n3165), .C(n3847), .D(n3848), .Z(n3845) );
  CANR2X1 U4924 ( .A(result_copy[9]), .B(n5189), .C(result_copy[10]), .D(n4483), .Z(n3825) );
  CANR4CX1 U4925 ( .A(n3823), .B(n3177), .C(n3827), .D(n3828), .Z(n3826) );
  CANR2X1 U4926 ( .A(n4469), .B(n5189), .C(result_copy[16]), .D(n4483), .Z(
        n3855) );
  COND3X1 U4927 ( .A(n3190), .B(n3165), .C(n3858), .D(n3859), .Z(n3856) );
  CANR2X1 U4928 ( .A(n5189), .B(n3377), .C(result_copy[12]), .D(n3753), .Z(
        n3834) );
  COND3X1 U4929 ( .A(n3193), .B(n3165), .C(n3837), .D(n3838), .Z(n3835) );
  COND3X1 U4930 ( .A(n329), .B(n3772), .C(n3811), .D(n3812), .Z(n1613) );
  CANR2X1 U4931 ( .A(result_copy[6]), .B(n5189), .C(result_copy[7]), .D(n3753), 
        .Z(n3812) );
  CEOX1 U4932 ( .A(n3808), .B(n3814), .Z(n3813) );
  COND3X1 U4933 ( .A(n332), .B(n3772), .C(n3792), .D(n3793), .Z(n1617) );
  CANR2X1 U4934 ( .A(result_copy[2]), .B(n5189), .C(result_copy[3]), .D(n3753), 
        .Z(n3793) );
  CEOX1 U4935 ( .A(n3795), .B(n3790), .Z(n3794) );
  COND3X1 U4936 ( .A(n4143), .B(n3248), .C(n4232), .D(n4233), .Z(n1511) );
  CND2X1 U4937 ( .A(result_not[43]), .B(n4168), .Z(n4232) );
  CANR2X1 U4938 ( .A(\intadd_1/SUM[10] ), .B(n4484), .C(n4177), .D(n3251), .Z(
        n4233) );
  COND3X1 U4939 ( .A(n4143), .B(n3243), .C(n4236), .D(n4237), .Z(n1509) );
  CND2X1 U4940 ( .A(result_not[45]), .B(n4168), .Z(n4236) );
  CANR2X1 U4941 ( .A(\intadd_1/SUM[12] ), .B(n4484), .C(n4177), .D(n3246), .Z(
        n4237) );
  COND3X1 U4942 ( .A(n3772), .B(n3368), .C(n3850), .D(n3851), .Z(n1605) );
  CANR2X1 U4943 ( .A(result_copy[14]), .B(n5189), .C(n4469), .D(n3753), .Z(
        n3851) );
  CENX1 U4944 ( .A(n3846), .B(n3853), .Z(n3852) );
  COND3X1 U4945 ( .A(n3772), .B(n3371), .C(n3839), .D(n3840), .Z(n1607) );
  CANR2X1 U4946 ( .A(result_copy[12]), .B(n5189), .C(result_copy[13]), .D(
        n4483), .Z(n3840) );
  CENX1 U4947 ( .A(n3842), .B(n3836), .Z(n3841) );
  COND3X1 U4948 ( .A(n3772), .B(n3372), .C(n3860), .D(n3861), .Z(n1603) );
  CANR2X1 U4949 ( .A(result_copy[16]), .B(n5189), .C(result_copy[17]), .D(
        n4483), .Z(n3861) );
  CENX1 U4950 ( .A(n3863), .B(n3857), .Z(n3862) );
  CANR11X1 U4951 ( .A(n3099), .B(n4921), .C(n3492), .D(n5192), .Z(n3594) );
  CANR11X1 U4952 ( .A(n3098), .B(n4928), .C(n3492), .D(n5192), .Z(n3584) );
  CANR11X1 U4953 ( .A(n3096), .B(n4875), .C(n3492), .D(n5192), .Z(n3564) );
  CANR11X1 U4954 ( .A(n3097), .B(n4863), .C(n3492), .D(n5192), .Z(n3574) );
  CANR11X1 U4955 ( .A(n3095), .B(n4868), .C(n3492), .D(n5192), .Z(n3554) );
  COND1XL U4956 ( .A(n3454), .B(n4477), .C(n3591), .Z(n235) );
  CANR4CX1 U4957 ( .A(n3592), .B(n3590), .C(n4895), .D(n3593), .Z(n3591) );
  CNR3XL U4958 ( .A(n4476), .B(n4921), .C(n3596), .Z(n3592) );
  CNR3XL U4959 ( .A(n3594), .B(n4895), .C(n3098), .Z(n3593) );
  CENX1 U4960 ( .A(n3136), .B(n4875), .Z(n3690) );
  COND2X1 U4961 ( .A(n4485), .B(n1741), .C(n3272), .D(n4482), .Z(n3973) );
  CND2X1 U4962 ( .A(n3738), .B(n3438), .Z(n3741) );
  COND4CX1 U4963 ( .A(n3738), .B(n3283), .C(n3740), .D(i[4]), .Z(n3742) );
  COND11X1 U4964 ( .A(n3360), .B(i[3]), .C(n3081), .D(n3739), .Z(n1652) );
  CND2X1 U4965 ( .A(i[3]), .B(n3740), .Z(n3739) );
  COND2X1 U4966 ( .A(n3647), .B(\intadd_0/B[10] ), .C(n4480), .D(n3678), .Z(
        n1675) );
  CENX1 U4967 ( .A(n3679), .B(n3120), .Z(n3678) );
  COND2X1 U4968 ( .A(n4481), .B(\intadd_0/B[14] ), .C(n4480), .D(n3689), .Z(
        n1671) );
  CENX1 U4969 ( .A(n3688), .B(n3690), .Z(n3689) );
  COND2X1 U4970 ( .A(n4481), .B(\intadd_0/B[18] ), .C(n4480), .D(n3700), .Z(
        n1667) );
  CENX1 U4971 ( .A(n3701), .B(n3114), .Z(n3700) );
  COND1XL U4972 ( .A(n4481), .B(\intadd_0/B[16] ), .C(n3694), .Z(n1669) );
  COND3X1 U4973 ( .A(n3116), .B(n3695), .C(n3696), .D(n3647), .Z(n3694) );
  COND1XL U4974 ( .A(n4481), .B(\intadd_0/B[12] ), .C(n3683), .Z(n1673) );
  COND3X1 U4975 ( .A(n3119), .B(n3684), .C(n3685), .D(n4481), .Z(n3683) );
  COND1XL U4976 ( .A(n4481), .B(\intadd_0/B[20] ), .C(n3705), .Z(n1665) );
  COND3X1 U4977 ( .A(n3113), .B(n3706), .C(n3707), .D(n4481), .Z(n3705) );
  CANR2X1 U4978 ( .A(n3817), .B(n3778), .C(n5180), .D(n5035), .Z(n3815) );
  CANR2X1 U4979 ( .A(result_copy[7]), .B(n5189), .C(n4483), .D(n3379), .Z(
        n3816) );
  CANR4CX1 U4980 ( .A(n3814), .B(n3808), .C(n3818), .D(n3819), .Z(n3817) );
  COND3X1 U4981 ( .A(n3772), .B(n3290), .C(n3796), .D(n3797), .Z(n1616) );
  CANR2X1 U4982 ( .A(result_copy[3]), .B(n5189), .C(n4483), .D(n3378), .Z(
        n3797) );
  CANR4CX1 U4983 ( .A(n3795), .B(n3790), .C(n3799), .D(n3800), .Z(n3798) );
  COND3X1 U4984 ( .A(n4143), .B(n3313), .C(n4212), .D(n4213), .Z(n1521) );
  CND2X1 U4985 ( .A(result_not[33]), .B(n4168), .Z(n4212) );
  CANR2X1 U4986 ( .A(\intadd_1/SUM[0] ), .B(n5177), .C(n4177), .D(n3316), .Z(
        n4213) );
  COND3X1 U4987 ( .A(n4143), .B(n3268), .C(n4216), .D(n4217), .Z(n1519) );
  CND2X1 U4988 ( .A(result_not[35]), .B(n4168), .Z(n4216) );
  CANR2X1 U4989 ( .A(\intadd_1/SUM[2] ), .B(n4484), .C(n4177), .D(n3272), .Z(
        n4217) );
  COND3X1 U4990 ( .A(n4143), .B(n3263), .C(n4220), .D(n4221), .Z(n1517) );
  CND2X1 U4991 ( .A(result_not[37]), .B(n4168), .Z(n4220) );
  CANR2X1 U4992 ( .A(\intadd_1/SUM[4] ), .B(n4484), .C(n4177), .D(n3266), .Z(
        n4221) );
  COND3X1 U4993 ( .A(n4143), .B(n3258), .C(n4224), .D(n4225), .Z(n1515) );
  CND2X1 U4994 ( .A(result_not[39]), .B(n4168), .Z(n4224) );
  CANR2X1 U4995 ( .A(\intadd_1/SUM[6] ), .B(n5177), .C(n4177), .D(n3261), .Z(
        n4225) );
  COND3X1 U4996 ( .A(n4143), .B(n3253), .C(n4228), .D(n4229), .Z(n1513) );
  CND2X1 U4997 ( .A(result_not[41]), .B(n4168), .Z(n4228) );
  CANR2X1 U4998 ( .A(\intadd_1/SUM[8] ), .B(n4484), .C(n4177), .D(n3256), .Z(
        n4229) );
  COND3X1 U4999 ( .A(n3772), .B(n3369), .C(n3892), .D(n3893), .Z(n1597) );
  CANR2X1 U5000 ( .A(result_copy[22]), .B(n5189), .C(result_copy[23]), .D(
        n4483), .Z(n3893) );
  CENX1 U5001 ( .A(n3888), .B(n3895), .Z(n3894) );
  COND3X1 U5002 ( .A(n3772), .B(n3374), .C(n3871), .D(n3872), .Z(n1601) );
  CANR2X1 U5003 ( .A(result_copy[18]), .B(n5189), .C(result_copy[19]), .D(
        n4483), .Z(n3872) );
  CENX1 U5004 ( .A(n3867), .B(n3874), .Z(n3873) );
  COND3X1 U5005 ( .A(n3772), .B(n3375), .C(n3881), .D(n3882), .Z(n1599) );
  CANR2X1 U5006 ( .A(result_copy[20]), .B(n5189), .C(result_copy[21]), .D(
        n4483), .Z(n3882) );
  CENX1 U5007 ( .A(n3884), .B(n3878), .Z(n3883) );
  COND3X1 U5008 ( .A(n3772), .B(n3481), .C(n3781), .D(n3782), .Z(n1619) );
  CANR2X1 U5009 ( .A(n5189), .B(n4488), .C(result_copy[1]), .D(n5191), .Z(
        n3782) );
  CANR1XL U5010 ( .A(n3785), .B(n3774), .C(n3786), .Z(n3784) );
  COND3X1 U5011 ( .A(n3772), .B(n3480), .C(n3801), .D(n3802), .Z(n1615) );
  CANR2X1 U5012 ( .A(n5189), .B(n3378), .C(result_copy[5]), .D(n5191), .Z(
        n3802) );
  CEOX1 U5013 ( .A(n3804), .B(n3800), .Z(n3803) );
  COND3X1 U5014 ( .A(n3772), .B(n3370), .C(n3820), .D(n3821), .Z(n1611) );
  CANR2X1 U5015 ( .A(n5189), .B(n3379), .C(result_copy[9]), .D(n5191), .Z(
        n3821) );
  CENX1 U5016 ( .A(n3823), .B(n3819), .Z(n3822) );
  COND4CX1 U5017 ( .A(n5192), .B(n3585), .C(n3589), .D(n3156), .Z(n3588) );
  COND4CX1 U5018 ( .A(n5192), .B(n3098), .C(n3590), .D(n4928), .Z(n3587) );
  CNR2X1 U5019 ( .A(n3585), .B(n3103), .Z(n3589) );
  COND4CX1 U5020 ( .A(n5192), .B(n3565), .C(n3569), .D(n3152), .Z(n3568) );
  COND4CX1 U5021 ( .A(n5192), .B(n3096), .C(n3570), .D(n4875), .Z(n3567) );
  CNR2X1 U5022 ( .A(n3565), .B(n3103), .Z(n3569) );
  COND3X1 U5023 ( .A(n4143), .B(n3247), .C(n4234), .D(n4235), .Z(n1510) );
  CND2X1 U5024 ( .A(result_not[44]), .B(n4168), .Z(n4234) );
  CANR2X1 U5025 ( .A(\intadd_1/SUM[11] ), .B(n4484), .C(n4177), .D(n3464), .Z(
        n4235) );
  COND3X1 U5026 ( .A(n4143), .B(n3252), .C(n4230), .D(n4231), .Z(n1512) );
  CND2X1 U5027 ( .A(result_not[42]), .B(n4168), .Z(n4230) );
  CANR2X1 U5028 ( .A(\intadd_1/SUM[9] ), .B(n5177), .C(n4177), .D(n3465), .Z(
        n4231) );
  COND3X1 U5029 ( .A(n4143), .B(n3257), .C(n4226), .D(n4227), .Z(n1514) );
  CND2X1 U5030 ( .A(result_not[40]), .B(n4168), .Z(n4226) );
  CANR2X1 U5031 ( .A(\intadd_1/SUM[7] ), .B(n3958), .C(n4177), .D(n3466), .Z(
        n4227) );
  COND3X1 U5032 ( .A(n3367), .B(n5184), .C(n4313), .D(n4314), .Z(n1478) );
  CND2X1 U5033 ( .A(result[12]), .B(n3078), .Z(n4314) );
  COND3X1 U5034 ( .A(result_not[12]), .B(n3353), .C(n4315), .D(n4475), .Z(
        n4313) );
  COND3X1 U5035 ( .A(n3371), .B(n5184), .C(n4319), .D(n4320), .Z(n1476) );
  CND2X1 U5036 ( .A(result[14]), .B(n3078), .Z(n4320) );
  COND3X1 U5037 ( .A(result_not[14]), .B(n3351), .C(n4321), .D(n5183), .Z(
        n4319) );
  COND3X1 U5038 ( .A(n3368), .B(n5184), .C(n4325), .D(n4326), .Z(n1474) );
  CND2X1 U5039 ( .A(result[16]), .B(n3078), .Z(n4326) );
  COND3X1 U5040 ( .A(result_not[16]), .B(n3349), .C(n4327), .D(n5183), .Z(
        n4325) );
  COND3X1 U5041 ( .A(n3372), .B(n4281), .C(n4331), .D(n4332), .Z(n1472) );
  CND2X1 U5042 ( .A(result[18]), .B(n3078), .Z(n4332) );
  COND3X1 U5043 ( .A(result_not[18]), .B(n3347), .C(n4333), .D(n5183), .Z(
        n4331) );
  COND3X1 U5044 ( .A(n3374), .B(n5184), .C(n4337), .D(n4338), .Z(n1470) );
  CND2X1 U5045 ( .A(result[20]), .B(n3078), .Z(n4338) );
  COND3X1 U5046 ( .A(result_not[20]), .B(n3345), .C(n4339), .D(n5183), .Z(
        n4337) );
  COND3X1 U5047 ( .A(n3288), .B(n5184), .C(n4316), .D(n4317), .Z(n1477) );
  CND2X1 U5048 ( .A(result[13]), .B(n3078), .Z(n4317) );
  COND3X1 U5049 ( .A(n3352), .B(result_not[13]), .C(n4318), .D(n4309), .Z(
        n4316) );
  COND3X1 U5050 ( .A(n3297), .B(n5184), .C(n4322), .D(n4323), .Z(n1475) );
  CND2X1 U5051 ( .A(result[15]), .B(n3078), .Z(n4323) );
  COND3X1 U5052 ( .A(n3350), .B(result_not[15]), .C(n4324), .D(n4475), .Z(
        n4322) );
  COND3X1 U5053 ( .A(n3287), .B(n5184), .C(n4328), .D(n4329), .Z(n1473) );
  CND2X1 U5054 ( .A(result[17]), .B(n3078), .Z(n4329) );
  COND3X1 U5055 ( .A(n3348), .B(result_not[17]), .C(n4330), .D(n5183), .Z(
        n4328) );
  COND3X1 U5056 ( .A(n3295), .B(n5184), .C(n4334), .D(n4335), .Z(n1471) );
  CND2X1 U5057 ( .A(result[19]), .B(n3078), .Z(n4335) );
  COND3X1 U5058 ( .A(n3346), .B(result_not[19]), .C(n4336), .D(n5183), .Z(
        n4334) );
  COND3X1 U5059 ( .A(n3772), .B(n3296), .C(n3885), .D(n3886), .Z(n1598) );
  CANR2X1 U5060 ( .A(result_copy[21]), .B(n5189), .C(result_copy[22]), .D(
        n4483), .Z(n3886) );
  COND3X1 U5061 ( .A(n3186), .B(n3165), .C(n3889), .D(n3890), .Z(n3887) );
  CANR2X1 U5062 ( .A(result_copy[19]), .B(n5189), .C(result_copy[20]), .D(
        n3753), .Z(n3876) );
  COND3X1 U5063 ( .A(n3187), .B(n3165), .C(n3879), .D(n3880), .Z(n3877) );
  COND3X1 U5064 ( .A(n3772), .B(n3295), .C(n3864), .D(n3865), .Z(n1602) );
  CANR2X1 U5065 ( .A(result_copy[17]), .B(n5189), .C(result_copy[18]), .D(
        n3753), .Z(n3865) );
  COND3X1 U5066 ( .A(n3189), .B(n3165), .C(n3868), .D(n3869), .Z(n3866) );
  CANR2X1 U5067 ( .A(result_copy[23]), .B(n5189), .C(result_copy[24]), .D(
        n4483), .Z(n3897) );
  COND3X1 U5068 ( .A(n3184), .B(n3165), .C(n3900), .D(n3901), .Z(n3898) );
  CND2X1 U5069 ( .A(n260), .B(n3414), .Z(n4150) );
  COND1XL U5070 ( .A(n3450), .B(n4477), .C(n3581), .Z(n237) );
  CANR1XL U5071 ( .A(n4899), .B(n3582), .C(n3583), .Z(n3581) );
  CNR3XL U5072 ( .A(n3584), .B(n4899), .C(n3097), .Z(n3583) );
  COND11X1 U5073 ( .A(n4476), .B(n4928), .C(n3585), .D(n3580), .Z(n3582) );
  COND1XL U5074 ( .A(n3448), .B(n4477), .C(n3561), .Z(n241) );
  CANR1XL U5075 ( .A(n4865), .B(n3562), .C(n3563), .Z(n3561) );
  CNR3XL U5076 ( .A(n3564), .B(n4865), .C(n3095), .Z(n3563) );
  COND11X1 U5077 ( .A(n4476), .B(n4875), .C(n3565), .D(n3560), .Z(n3562) );
  COND1XL U5078 ( .A(n3442), .B(n4477), .C(n3571), .Z(n239) );
  CANR4CX1 U5079 ( .A(n3572), .B(n3570), .C(n4836), .D(n3573), .Z(n3571) );
  CNR3XL U5080 ( .A(n4476), .B(n4863), .C(n3576), .Z(n3572) );
  CNR3XL U5081 ( .A(n3574), .B(n4836), .C(n3096), .Z(n3573) );
  COND1XL U5082 ( .A(n3735), .B(n3440), .C(n3748), .Z(n1624) );
  CANR11X1 U5083 ( .A(n3738), .B(n3440), .C(i[0]), .D(n3083), .Z(n3748) );
  COND4CX1 U5084 ( .A(n3735), .B(n3736), .C(n3437), .D(n3737), .Z(n1653) );
  CND2X1 U5085 ( .A(n3738), .B(n3440), .Z(n3736) );
  CND2X1 U5086 ( .A(\cust[1] ), .B(n284), .Z(n3752) );
  CENX1 U5087 ( .A(n5141), .B(n4479), .Z(n4090) );
  CENX1 U5088 ( .A(opera2[55]), .B(n4478), .Z(n4103) );
  CENX1 U5089 ( .A(opera2[59]), .B(n4478), .Z(n4129) );
  CANR3X1 U5090 ( .A(\cust[1] ), .B(n3479), .C(n4173), .D(n4165), .Z(n4172) );
  CNR3XL U5091 ( .A(n3389), .B(n3475), .C(n4170), .Z(n4173) );
  COND3X1 U5092 ( .A(n4143), .B(n3267), .C(n4218), .D(n4219), .Z(n1518) );
  CND2X1 U5093 ( .A(result_not[36]), .B(n4168), .Z(n4218) );
  CANR2X1 U5094 ( .A(\intadd_1/SUM[3] ), .B(n4484), .C(n1741), .D(n4177), .Z(
        n4219) );
  CANR11X1 U5095 ( .A(n3126), .B(n4977), .C(n3492), .D(n5192), .Z(n3624) );
  CANR11X1 U5096 ( .A(n3635), .B(n4971), .C(n3492), .D(n5192), .Z(n3634) );
  CANR11X1 U5097 ( .A(n3101), .B(n4923), .C(n3492), .D(n5192), .Z(n3604) );
  CANR11X1 U5098 ( .A(n3102), .B(n4969), .C(n3492), .D(n5192), .Z(n3614) );
  CEOX1 U5099 ( .A(n3482), .B(opera1_copy[0]), .Z(n3945) );
  CENX1 U5100 ( .A(n3136), .B(n4818), .Z(n3712) );
  COND1XL U5101 ( .A(n3467), .B(n4477), .C(n3631), .Z(n227) );
  CANR4CX1 U5102 ( .A(n3632), .B(n3630), .C(n4943), .D(n3633), .Z(n3631) );
  CNR3XL U5103 ( .A(n4476), .B(n4971), .C(n3131), .Z(n3632) );
  CNR3XL U5104 ( .A(n3634), .B(n4943), .C(n3126), .Z(n3633) );
  CNR2X1 U5105 ( .A(n4480), .B(n4986), .Z(n3488) );
  COND11X1 U5106 ( .A(n4167), .B(n4477), .C(n4166), .D(n4168), .Z(n1557) );
  COND1XL U5107 ( .A(n3394), .B(n4150), .C(valid), .Z(n4167) );
  COND1XL U5108 ( .A(n3462), .B(n4477), .C(n3601), .Z(n233) );
  CANR1XL U5109 ( .A(n4920), .B(n3602), .C(n3603), .Z(n3601) );
  CNR3XL U5110 ( .A(n3604), .B(n4920), .C(n3099), .Z(n3603) );
  COND11X1 U5111 ( .A(n4476), .B(n4923), .C(n3605), .D(n3600), .Z(n3602) );
  COND2X1 U5112 ( .A(n3165), .B(n3197), .C(n3178), .D(n4524), .Z(n3791) );
  COND2X1 U5113 ( .A(n3647), .B(\intadd_0/B[2] ), .C(n4480), .D(n3656), .Z(
        n1683) );
  CENX1 U5114 ( .A(n3657), .B(n3129), .Z(n3656) );
  COND2X1 U5115 ( .A(n3647), .B(\intadd_0/B[0] ), .C(n4480), .D(n3651), .Z(
        n1685) );
  CENX1 U5116 ( .A(n3650), .B(n3652), .Z(n3651) );
  COND2X1 U5117 ( .A(n4481), .B(\intadd_0/B[6] ), .C(n4480), .D(n3667), .Z(
        n1679) );
  CENX1 U5118 ( .A(n3666), .B(n3668), .Z(n3667) );
  COND1XL U5119 ( .A(n4481), .B(\intadd_0/B[8] ), .C(n3672), .Z(n1677) );
  COND3X1 U5120 ( .A(n3122), .B(n3673), .C(n3674), .D(n4481), .Z(n3672) );
  CND3XL U5121 ( .A(n284), .B(n4793), .C(n3751), .Z(n3754) );
  CNIVX1 U5122 ( .A(n3776), .Z(n5180) );
  CNR3XL U5123 ( .A(muordi), .B(n4479), .C(n4476), .Z(n3776) );
  CND3XL U5124 ( .A(n3492), .B(cin1a), .C(n3644), .Z(n3642) );
  COND4CX1 U5125 ( .A(n5192), .B(n3635), .C(n3640), .D(n4971), .Z(n3637) );
  COND4CX1 U5126 ( .A(n5192), .B(n3131), .C(n3639), .D(n3164), .Z(n3638) );
  CNR2X1 U5127 ( .A(n3131), .B(n3103), .Z(n3639) );
  COND4CX1 U5128 ( .A(n5192), .B(n3625), .C(n3629), .D(n3162), .Z(n3628) );
  COND4CX1 U5129 ( .A(n5192), .B(n3126), .C(n3630), .D(n4977), .Z(n3627) );
  CNR2X1 U5130 ( .A(n3625), .B(n3103), .Z(n3629) );
  COND4CX1 U5131 ( .A(n5192), .B(n3605), .C(n3609), .D(n3159), .Z(n3608) );
  COND4CX1 U5132 ( .A(n5192), .B(n3101), .C(n3610), .D(n4923), .Z(n3607) );
  CNR2X1 U5133 ( .A(n3605), .B(n3103), .Z(n3609) );
  COND3X1 U5134 ( .A(n3370), .B(n5184), .C(n4306), .D(n4307), .Z(n1480) );
  CND2X1 U5135 ( .A(result[10]), .B(n3078), .Z(n4307) );
  COND3X1 U5136 ( .A(result_not[10]), .B(n3355), .C(n4308), .D(n4475), .Z(
        n4306) );
  COND3X1 U5137 ( .A(n327), .B(n5184), .C(n4310), .D(n4311), .Z(n1479) );
  CND2X1 U5138 ( .A(result[11]), .B(n3078), .Z(n4311) );
  COND3X1 U5139 ( .A(n3354), .B(result_not[11]), .C(n4312), .D(n5183), .Z(
        n4310) );
  COND2X1 U5140 ( .A(n3365), .B(n4281), .C(n4474), .D(n4299), .Z(n4298) );
  COND4CX1 U5141 ( .A(n3357), .B(result_not[6]), .C(result_not[7]), .D(n4300), 
        .Z(n4299) );
  COND2X1 U5142 ( .A(n3289), .B(n4281), .C(n4474), .D(n4304), .Z(n4303) );
  COND4CX1 U5143 ( .A(n3356), .B(result_not[8]), .C(result_not[9]), .D(n4305), 
        .Z(n4304) );
  COND1XL U5144 ( .A(n4481), .B(\intadd_0/B[4] ), .C(n3661), .Z(n1681) );
  COND3X1 U5145 ( .A(n3125), .B(n3662), .C(n3663), .D(n4481), .Z(n3661) );
  COND1XL U5146 ( .A(result_copy[1]), .B(n5185), .C(n4178), .Z(n1553) );
  CANR2X1 U5147 ( .A(result_not[1]), .B(n4168), .C(n4179), .D(n335), .Z(n4178)
         );
  COND1XL U5148 ( .A(result_copy[3]), .B(n5185), .C(n4181), .Z(n1551) );
  CANR2X1 U5149 ( .A(result_not[3]), .B(n4168), .C(n4179), .D(n3481), .Z(n4181) );
  COND1XL U5150 ( .A(result_copy[5]), .B(n5185), .C(n4183), .Z(n1549) );
  COND1XL U5151 ( .A(result_copy[7]), .B(n5185), .C(n4185), .Z(n1547) );
  CANR2X1 U5152 ( .A(result_not[7]), .B(n4168), .C(n4179), .D(n3480), .Z(n4185) );
  COND1XL U5153 ( .A(result_copy[9]), .B(n5185), .C(n4187), .Z(n1545) );
  COND1XL U5154 ( .A(n5185), .B(n3377), .C(n4189), .Z(n1543) );
  CANR2X1 U5155 ( .A(result_not[11]), .B(n4168), .C(n4179), .D(n3370), .Z(
        n4189) );
  COND1XL U5156 ( .A(result_copy[13]), .B(n5185), .C(n4191), .Z(n1541) );
  CANR2X1 U5157 ( .A(result_not[13]), .B(n5186), .C(n4179), .D(n3367), .Z(
        n4191) );
  COND1XL U5158 ( .A(n4469), .B(n5185), .C(n4193), .Z(n1539) );
  CANR2X1 U5159 ( .A(result_not[15]), .B(n5186), .C(n4179), .D(n3371), .Z(
        n4193) );
  COND1XL U5160 ( .A(result_copy[17]), .B(n5185), .C(n4195), .Z(n1537) );
  CANR2X1 U5161 ( .A(result_not[17]), .B(n5186), .C(n4179), .D(n3368), .Z(
        n4195) );
  COND1XL U5162 ( .A(result_copy[19]), .B(n5185), .C(n4197), .Z(n1535) );
  CANR2X1 U5163 ( .A(result_not[19]), .B(n5186), .C(n4179), .D(n3372), .Z(
        n4197) );
  COND1XL U5164 ( .A(result_copy[21]), .B(n5185), .C(n4199), .Z(n1533) );
  CANR2X1 U5165 ( .A(result_not[21]), .B(n5186), .C(n4179), .D(n3374), .Z(
        n4199) );
  COND1XL U5166 ( .A(result_copy[23]), .B(n5185), .C(n4201), .Z(n1531) );
  CANR2X1 U5167 ( .A(result_not[23]), .B(n5186), .C(n4179), .D(n3375), .Z(
        n4201) );
  COND1XL U5168 ( .A(result_copy[25]), .B(n5185), .C(n4203), .Z(n1529) );
  CANR2X1 U5169 ( .A(result_not[25]), .B(n5186), .C(n4179), .D(n3369), .Z(
        n4203) );
  COND1XL U5170 ( .A(result_copy[27]), .B(n5185), .C(n4205), .Z(n1527) );
  CANR2X1 U5171 ( .A(result_not[27]), .B(n5186), .C(n4179), .D(n3366), .Z(
        n4205) );
  COND1XL U5172 ( .A(result_copy[29]), .B(n5185), .C(n4207), .Z(n1525) );
  CANR2X1 U5173 ( .A(result_not[29]), .B(n5186), .C(n4179), .D(n3376), .Z(
        n4207) );
  COND1XL U5174 ( .A(n5009), .B(n5185), .C(n4209), .Z(n1523) );
  CANR2X1 U5175 ( .A(result_not[31]), .B(n5186), .C(n4179), .D(n3373), .Z(
        n4209) );
  COND1XL U5176 ( .A(n4481), .B(n3474), .C(n3649), .Z(n1686) );
  COND3X1 U5177 ( .A(cin1b), .B(n3644), .C(n3650), .D(n4481), .Z(n3649) );
  COND1XL U5178 ( .A(n3471), .B(n4477), .C(n4950), .Z(n229) );
  CANR1XL U5179 ( .A(n4952), .B(n3622), .C(n3623), .Z(n3621) );
  COND11X1 U5180 ( .A(n4476), .B(n4977), .C(n3625), .D(n3620), .Z(n3622) );
  CNR3XL U5181 ( .A(n3624), .B(n4952), .C(n3102), .Z(n3623) );
  COND1XL U5182 ( .A(result_copy[2]), .B(n5185), .C(n4180), .Z(n1552) );
  CANR2X1 U5183 ( .A(result_not[2]), .B(n4168), .C(n4179), .D(n3291), .Z(n4180) );
  COND1XL U5184 ( .A(n5185), .B(n3378), .C(n4182), .Z(n1550) );
  CANR2X1 U5185 ( .A(result_not[4]), .B(n4168), .C(n4179), .D(n3364), .Z(n4182) );
  COND1XL U5186 ( .A(result_copy[6]), .B(n5185), .C(n4184), .Z(n1548) );
  CANR2X1 U5187 ( .A(result_not[6]), .B(n4168), .C(n4179), .D(n3290), .Z(n4184) );
  COND1XL U5188 ( .A(n5185), .B(n3379), .C(n4186), .Z(n1546) );
  CANR2X1 U5189 ( .A(result_not[8]), .B(n4168), .C(n4179), .D(n3365), .Z(n4186) );
  COND1XL U5190 ( .A(result_copy[10]), .B(n5185), .C(n4188), .Z(n1544) );
  CANR2X1 U5191 ( .A(result_not[10]), .B(n4168), .C(n4179), .D(n3289), .Z(
        n4188) );
  COND1XL U5192 ( .A(result_copy[12]), .B(n5185), .C(n4190), .Z(n1542) );
  CANR2X1 U5193 ( .A(result_not[12]), .B(n5186), .C(n327), .D(n4179), .Z(n4190) );
  COND1XL U5194 ( .A(result_copy[14]), .B(n5185), .C(n4192), .Z(n1540) );
  CANR2X1 U5195 ( .A(result_not[14]), .B(n5186), .C(n4179), .D(n3288), .Z(
        n4192) );
  COND1XL U5196 ( .A(n3455), .B(n4477), .C(n3611), .Z(n231) );
  CANR4CX1 U5197 ( .A(n3612), .B(n3610), .C(n4935), .D(n3613), .Z(n3611) );
  CNR3XL U5198 ( .A(n4476), .B(n4969), .C(n3616), .Z(n3612) );
  CNR3XL U5199 ( .A(n3614), .B(n4935), .C(n3101), .Z(n3613) );
  COND1XL U5200 ( .A(result_copy[16]), .B(n5185), .C(n4194), .Z(n1538) );
  CANR2X1 U5201 ( .A(result_not[16]), .B(n5186), .C(n4179), .D(n3297), .Z(
        n4194) );
  COND1XL U5202 ( .A(result_copy[18]), .B(n5185), .C(n4196), .Z(n1536) );
  CANR2X1 U5203 ( .A(result_not[18]), .B(n5186), .C(n4179), .D(n3287), .Z(
        n4196) );
  COND1XL U5204 ( .A(result_copy[20]), .B(n5185), .C(n4198), .Z(n1534) );
  CANR2X1 U5205 ( .A(result_not[20]), .B(n5186), .C(n4179), .D(n3295), .Z(
        n4198) );
  COND1XL U5206 ( .A(result_copy[22]), .B(n5185), .C(n4200), .Z(n1532) );
  CANR2X1 U5207 ( .A(result_not[22]), .B(n5186), .C(n4179), .D(n3294), .Z(
        n4200) );
  COND1XL U5208 ( .A(result_copy[24]), .B(n5185), .C(n4202), .Z(n1530) );
  CANR2X1 U5209 ( .A(result_not[24]), .B(n5186), .C(n4179), .D(n3296), .Z(
        n4202) );
  COND1XL U5210 ( .A(result_copy[26]), .B(n5185), .C(n4204), .Z(n1528) );
  CANR2X1 U5211 ( .A(result_not[26]), .B(n5186), .C(n4179), .D(n3286), .Z(
        n4204) );
  COND1XL U5212 ( .A(result_copy[28]), .B(n5185), .C(n4206), .Z(n1526) );
  CANR2X1 U5213 ( .A(result_not[28]), .B(n5186), .C(n4179), .D(n3285), .Z(
        n4206) );
  COND1XL U5214 ( .A(result_copy[30]), .B(n5185), .C(n4208), .Z(n1524) );
  CANR2X1 U5215 ( .A(result_not[30]), .B(n5186), .C(n4179), .D(n3293), .Z(
        n4208) );
  COND1XL U5216 ( .A(n3080), .B(n3363), .C(n3646), .Z(n1687) );
  CANR1XL U5217 ( .A(n3415), .B(n3080), .C(n4481), .Z(n3646) );
  COND4CX1 U5218 ( .A(n4170), .B(n4168), .C(n3648), .D(n4171), .Z(n1555) );
  CND2X1 U5219 ( .A(n3648), .B(n5005), .Z(n4171) );
  CAN2X1 U5220 ( .A(n4179), .B(n1770), .Z(n3958) );
  CAN2X1 U5221 ( .A(n4179), .B(n1770), .Z(n5177) );
  COND4CX1 U5222 ( .A(n3774), .B(n3775), .C(n5180), .D(n4708), .Z(n3773) );
  COND2X1 U5223 ( .A(n332), .B(n4281), .C(n4292), .D(n4474), .Z(n4291) );
  CENX1 U5224 ( .A(n3358), .B(result_not[4]), .Z(n4292) );
  COND2X1 U5225 ( .A(n329), .B(n4281), .C(n4302), .D(n4474), .Z(n4301) );
  CENX1 U5226 ( .A(n3356), .B(result_not[8]), .Z(n4302) );
  COND2X1 U5227 ( .A(n335), .B(n4281), .C(n4282), .D(n4474), .Z(n4280) );
  CENX1 U5228 ( .A(result_not[0]), .B(cina), .Z(n4282) );
  COND2X1 U5229 ( .A(n3481), .B(n4281), .C(n4287), .D(n4474), .Z(n4286) );
  CENX1 U5230 ( .A(result_not[2]), .B(n3359), .Z(n4287) );
  COND2X1 U5231 ( .A(n3480), .B(n4281), .C(n4297), .D(n4474), .Z(n4296) );
  CENX1 U5232 ( .A(result_not[6]), .B(n3357), .Z(n4297) );
  COND2X1 U5233 ( .A(n3291), .B(n4281), .C(n4474), .D(n4284), .Z(n4283) );
  COND4CX1 U5234 ( .A(cina), .B(result_not[0]), .C(result_not[1]), .D(n4285), 
        .Z(n4284) );
  COND2X1 U5235 ( .A(n3364), .B(n4281), .C(n4474), .D(n4289), .Z(n4288) );
  COND4CX1 U5236 ( .A(n3359), .B(result_not[2]), .C(result_not[3]), .D(n4290), 
        .Z(n4289) );
  COND2X1 U5237 ( .A(n3290), .B(n4281), .C(n4474), .D(n4294), .Z(n4293) );
  COND4CX1 U5238 ( .A(n3358), .B(result_not[4]), .C(result_not[5]), .D(n4295), 
        .Z(n4294) );
  CANR3X1 U5239 ( .A(n3648), .B(n4828), .C(n4165), .D(n4477), .Z(n4169) );
  CENX1 U5240 ( .A(n3136), .B(n4690), .Z(n3732) );
  CENX1 U5241 ( .A(n4478), .B(n5040), .Z(n3804) );
  CENX1 U5242 ( .A(n4478), .B(n5096), .Z(n3926) );
  CNR2X1 U5243 ( .A(n5008), .B(n5007), .Z(n259) );
  CNR2IX1 U5244 ( .B(n4828), .A(n5008), .Z(N145) );
  CIVXL U5245 ( .A(n4474), .Z(n5183) );
  CIVX1 U5246 ( .A(n4177), .Z(n5185) );
  CIVX2 U5247 ( .A(n4143), .Z(n5187) );
  CIVXL U5248 ( .A(n4485), .Z(n5188) );
  CIVXL U5249 ( .A(n4487), .Z(n5190) );
  CIVXL U5250 ( .A(n4482), .Z(n5191) );
endmodule

